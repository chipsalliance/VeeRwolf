0102829300000297
2840106F30529073
00112023FB010113
0041242300312223
0061282300512623
01C12C2300712A23
03E1202301D12E23
02A1242303F12223
02C1282302B12623
02E12C2302D12A23
0501202302F12E23
341022F305112223
300022F304512423
1BC000EF04512623
02051E6300000313
800003B7342022F3
0072F2B3FFF38393
00628A6300B00313
0000009700010513
1B00106F12408093
0042829304812283
0800006F04512423
0000339700010293
0043A1039D838393
00512023FF010113
001E0E130003AE03
3420257301C3A023
FFF28293800002B7
134000EF00557533
4342829300002297
00A282B300351513
0042A3030002A503
00003317000300E7
0003238398830313
00732023FFF38393
0002811300012283
02032E0300832383
00003297087E0863
0082A30396028293
0293282302832623
03332C2303232A23
0553202303432E23
0573242305632223
0593282305832623
05B32C2305A32A23
0000239702232423
0003AE037C438393
0202A30307C32623
028321030062A423
0303248302C32403
0383298303432903
04032A8303C32A03
04832B8304432B03
05032C8304C32C03
05832D8305432D03
3412907304812283
3002907304C12283
0041218300012083
00C1228300812203
0141238301012303
01C12E8301812E03
02412F8302012F03
02C1258302812503
0341268303012603
03C1278303812703
0441288304012803
3020007305010113
00A312B300100313
000080673442B373
80000337342022F3
000005130062F2B3
0015051300028463
0000007300008067
8442829300003297
06C323830082A303
300522F300857513
0000806700038513
0200079302060063
00F04C6340C787B3
00000713FE060513
0007059300A5D533
00C5D73300008067
00F595B300C55533
FE9FF06F00B56533
0006081300058793
0005031300068713
000028B728069663
0EC5F66375888893
0CE6786300010737
00C6B6B30FF00693
00D6573300369693
0008C70300E888B3
0200071300D706B3
00070C6340D70733
00D556B300E797B3
00F6E5B300E61833
0108551300E51333
0108161302A5F733
0103569301065613
0107171302A5D5B3
02B607B300D766B3
00F6FE6300058713
FFF58713010686B3
00F6F6630106E863
010686B3FFE58713
02A6F7B340F686B3
0103531301031313
0107979302A6D6B3
02D605B30067E333
00B37C6300068513
FFF6851300680333
00B3746301036663
01071713FFE68513
0000059300A76733
010007370E40006F
F2E66CE301000693
F31FF06F01800693
0010069300061663
000106B702C6D833
0FF006930CD87263
008007130106F463
00D888B300E856B3
00E686B30008C683
40D7073302000713
410787B30A071863
0108561300100593
0108D89301081893
02C7F73301035693
0107171302C7D7B3
02F8853300D766B3
00A6FE6300078713
FFF78713010686B3
00A6F6630106E863
010686B3FFE78713
02C6F7B340A686B3
0103531301031313
0107979302C6D6B3
02D888B30067E333
01137C6300068513
FFF6851300680333
0113746301036663
01071713FFE68513
0007051300A76733
010006B700008067
F4D862E301000713
F3DFF06F01800713
00D7D5B300E81833
00D556B300E51333
00E797B301085513
00F6E8B302A5F733
0107D79301081793
02A5D5B30108D613
00C7673301071713
0005861302B786B3
0107073300D77E63
01076863FFF58613
FFE5861300D77663
40D706B301070733
0108989302A6F733
02A6D6B30108D893
02D785B301071713
00068713011767B3
010787B300B7FE63
0107E863FFF68713
FFE6871300B7F663
40B787B3010787B3
00E5E5B301061593
18D5E663EB5FF06F
04E6F46300010737
00D835B30FF00813
0000273700359593
7587071300B6D833
0007480301070733
0200059300B80833
02059663410585B3
EEF6ECE300100713
0016471300C53633
01000737EEDFF06F
FCE6E0E301000593
FB9FF06F01800593
00B696B301065733
0106DE9300D766B3
03D778B30107D733
0105583300B797B3
0106979300F86333
010358130107D793
03D7573300B61633
0108E83301089893
00070E1302E78F33
00D8083301E87E63
00D86863FFF70E13
FFE70E1301E87663
41E8083300D80833
03D8583303D878B3
03078EB301089893
0107D79301031793
0008071300F8E7B3
00D787B301D7FE63
00D7E863FFF80713
FFE8071301D7F663
010E1E1300D787B3
00010EB741D787B3
FFFE881300EE6733
0107589301077333
0106561301067833
0308883303030E33
02C30333010E5693
006686B301030333
0106F46302C888B3
0106D61301D888B3
0317E663011608B3
000107B7CF179AE3
00F6F6B3FFF78793
00FE7E3301069693
01C686B300B51533
DAD57CE300000593
CC9FF06FFFF70713
0000071300000593
000035B7DA5FF06F
8585859300003537
7580006F86850513
0085530300452883
00A54F0300052803
FFF0079303130E33
0008859300F505A3
00C00F9300000613
01C8083302000E93
0000061301E64A63
0466CA6300000693
02BE57B300008067
03F6073300C52683
0047069300E68733
00D7242300D72223
00C505A300FEEC63
FFC5F5930025D593
FBDFF06F00160613
03D7C7B301F78793
0027979301072023
FDDFF06F00F80833
0005278300C52703
0047059300168693
00B7A02300C787B3
0116063300872583
0087258300B7A223
00F7242300F5A023
FF010113F7DFF06F
0005851300050793
0006861300060593
000780E700112623
0D9010EF674010EF
0000806700000513
00812423FF010113
0450051300050413
0091222300112623
000400E700058493
0520051300048593
00040313000400E7
00C1208300812403
0041248300048593
0101011305200513
0005A78300030067
00F5A02300178793
91C7A303000037B7
FB01011300030067
03312E2304812423
03512A2303412C23
0411262303712623
0521202304912223
0381242303612823
03A1202303912223
00050A1301B12E23
0006099300058A93
0010041300068B93
0007041300E05463
02000C1300100793
03000C1300FB9463
001009133B9AD4B7
0000079300A00B13
00100C93A0048493
00A00D1300200D93
0899E06300079463
000A85930299D533
0305051300190913
00100793000A00E7
0299F9B3FFFB0B13
FD9B1AE303A4D4B3
03098513000A8593
00300793000A00E7
06FB8A6341240433
0481240304C12083
0401290304412483
03812A0303C12983
03012B0303412A83
02812C0302C12B83
02012D0302412C83
0501011301C12D83
F9644EE300008067
000A8593F97DECE3
00F12623000C0513
00190913000A00E7
F7DFF06F00C12783
02000513000A8593
FFF40413000A00E7
F8DFF06FFE8048E3
90A7AE23000037B7
FB01011300008067
0491222304812423
03312E2305212023
03512A2303412C23
01B12E2303A12023
0361282304112623
0381242303712623
0005041303912223
00060A9300058493
0000091300068D93
00000A13FFF00993
000AC50300000D13
04C1208304051063
0441248304812403
03C1298304012903
03412A8303812A03
02C12B8303012B03
02412C8302812C03
01C12D8302012D03
0000806705010113
02500693000D1E63
000485933AD50863
001A8A93000400E7
06400693FA5FF06F
06A6E26312D50E63
02A6EA6303900693
0ED57C6303100693
38D5086302D00693
0CF5086303000793
02E5126302500713
0250051300048593
18C0006F000400E7
1ED5066305800693
32E50A6306300713
0250051300048593
00048593000400E7
FD5FF06F000AC503
1AD5026307000693
0690069302A6E863
06C006930CD50263
0680069300D50663
06800693FCD514E3
08A91E6308D51A63
F59FF06F04800913
12D5066307500693
0730071302A6EE63
000DAC03FAE510E3
000C0B13004D8B93
28051C63000B4503
00FA186300300793
41698B33418B0B33
000B8D9329604A63
078006930E80006F
07A0069314D50463
0009DE63F99FF06F
FD0509932A0A0E63
00200A13EE0A1AE3
FE09C8E3EEDFF06F
02D989B300A00693
013509B3FD098993
06C00693FE1FF06F
28A9086300D51463
00050913F20910E3
07A00713EBDFF06F
000DA60304E91263
02065063004D8D93
02D0051300048593
000400E700C12423
FFF9899300812603
0009871340C00633
00048593000A0693
C79FF0EF00040513
06C007130480006F
04C00713FAE90EE3
007D8793FAE91AE3
00072603FF87F713
00870D9300472683
00E6073380000737
00D7073300C73733
00048593F8070AE3
BCDFF0EF00040513
E29FF06F00000D13
00E9186307A00713
004D8D93000DA603
06C00713F8DFF06F
04C00713FEE908E3
007D8793FEE914E3
00870D93FF87F713
0047270300072603
FB1FF06FF60702E3
0300051300048593
00048593000400E7
000400E707800513
00100A1300800993
07000693000AC603
000DAB8300D61A63
004D8D9300000C13
06C006930280006F
04C00693FED906E3
007D8793FED912E3
0006AB83FF87F693
00868D930046AC03
00000C9301000793
04000B1300012423
000B0613FFCB0B13
000C0593000B8513
D8CFF0EF00F12623
00C1278300F57513
0081270306051663
0007146303000693
00A68533060B1863
0004859301851513
00F1242341855513
001C8C93000400E7
020B186300812783
00000D1300300693
00199713D0DA1AE3
ED905EE341970CB3
0200051300048593
FFFC8C93000400E7
01A12423FEDFF06F
00900713F79FF06F
FAA760E305700693
F99FF06F03000693
00E12623FFF78713
0010079300F9CC63
0004859300FA1C63
000400E703000513
F3DFF06F00C12783
FEFA1AE300200793
0200051300048593
00048593FE5FF06F
000400E7001B0B13
00048593D59FF06F
000400E702000513
D5DFF06FFFFB0B13
004D8B13000DA503
000400E700048593
E35FF06F000B0D93
FFF0099300000913
00100D1300000A13
00300A13C4DFF06F
00100A13C45FF06F
04C00913C3DFF06F
FE010113C35FF06F
0000153700050613
8245051300058693
00112E2300C10593
B61FF0EF00012623
0201011301C12083
FC01011300008067
0241059302B12223
02C1242300112E23
02E1282302D12623
03012C2302F12A23
00B1262303112E23
01C12083FA5FF0EF
0000806704010113
0080079300008067
304050733007B7F3
0000806734405073
00812423FF010113
0000343700912223
00A0079300112623
9984041300050493
0004250300F51C63
00D0059300452783
000780E70047A783
0045278300042503
0047A7830FF4F593
00C12083000780E7
0004851300812403
0101011300412483
FF01011300008067
0000143700812423
00112623E9040513
E904051350C000EF
00C1208300812403
A65FF06F01010113
00112623FF010113
87C5051300003537
000037B76A0000EF
FB9FF0EF98A7AC23
0000051300C12083
0000806701010113
0007A023F00C37B7
00478713F00C27B7
0007202312C78793
FEF71CE300470713
00478713F00C07B7
12C7879300F00693
0047071300D72023
F00C47B7FEF71CE3
12C7879300478713
0047071300072023
F00C57B7FEF71CE3
12C7879300478713
0047071300072023
BC905073FEF71CE3
BCC05073BCB05073
80078793000017B7
000005133047A7F3
FF01011300008067
0081242300112623
FC802473BCA05073
0FF4741300245413
9887AE23000037B7
03E00793FFF40713
0000051300E7F663
00B40713254000EF
00371713000027B7
00E787B351C78793
000706630047A703
000700E70007A503
40B78793000017B7
0024141300F40433
00F40433F00C07B7
00C1208300042023
0101011300812403
FF55071300008067
02E7E66303F00793
3007B7F300800793
F00C07377F550513
00E5053300251513
00E5202300100713
3007A7F30087F793
00B0071300008067
00A7746300050793
00100513FBDFF06F
3045257300F51533
800017B700008067
0207A5030247A703
FEE59AE30247A583
FE01011300008067
00112E2301212823
00912A2300812C23
0141242301312623
0080091301512223
00003A3730093973
FB9FF0EF988A0A13
004A2A83000A2403
4085053300050993
0005849300A9B7B3
415585B30007A637
0000069312060613
96CFF0EF40F585B3
120787930007A7B7
0089791302F50533
00F707B300850733
015506B300A73533
00D6063300E7B633
0137B5B3413789B3
00EA2023409604B3
40B484B300DA2223
0004966302904263
0135EC633E700593
24078793000F47B7
00E7B73300F707B3
8000173700D70633
02D72623FFF00693
02C7262302F72423
0181240330092973
0141248301C12083
00C1298301012903
00412A8300812A03
0201011300100513
FF01011319C0106F
ED9FF0EF00112623
120787930007A7B7
00F507B380001737
02D72623FFF00693
00B5053300A7B533
02A7262302F72423
E89FF0EF00700513
0000051300C12083
0000806701010113
0000051300008067
0080079300008067
000080673007A7F3
00112623FF010113
FF01011343C000EF
0005059300112623
00000513342027F3
FF010113424000EF
342027F300112623
0010051300000593
FF010113FC9FF0EF
444000EF00112623
4B8000EFBF5FF0EF
00050663F1402573
FFDFF06F10500073
E201011300002117
80028293000012B7
FC9FF0EF00510133
FD010113CF4FF06F
0007099301312E23
01412C2303012703
0008869300068A13
0291222302812423
0211262303212023
0005091300058413
00F1262300060493
3E9000EF01012423
FB04859300C12783
FF05F59300B405B3
000027B702F5A823
8807879300812803
000017B704F5A623
0281240302C12083
0345A4232B878793
0305AA230335A623
02B9242304F5A423
0201290302412483
01812A0301C12983
0000806703010113
0005C70300054783
0007966300E79463
0000806740E78533
0015859300150513
0FF5F693FE1FF06F
0037F71300050793
0FF5F59304071863
00B765B300859713
00B765B301059713
0007871300C78333
40E308B300300813
0026571303186E63
00B787B300271593
02B70733FFC00593
00E7873300C70733
0000806702E79463
00178793FE060EE3
FFF60613FED78FA3
00470713F9DFF06F
FB9FF06FFEB72E23
FED78FA300178793
FFF00513FD1FF06F
000037B700008067
0000806792A7A023
0080071300852803
0048268330073773
0606886300877713
0087A78300052783
060600630007A603
00C787B300369793
0085288302D7D7B3
00C5C6030008A583
080663130FF67613
0085230300658623
0047D59300032303
00B300230FF5F593
00C7D79300852583
0005A5830FF7F793
0085278300F58223
00C786230007A783
0085278300D8A223
0007A78300300693
0088478300D78623
0017F79300B00693
02B0069300078463
0007A78300852783
0085278300D78823
0007A783F8700693
0085278300D78423
0007C6830007A783
3007277300078223
0000806700000513
0007A70300852783
0017F79301474783
0007478300078A63
00F5802300000513
FFF0051300008067
0085278300008067
014706930007A703
0207F7930006C783
00B70023FE078CE3
0085278300008067
0147C5030007A783
00F5751300155513
0025171300008067
00150513000037B7
002515138A478793
00E78733FF010113
0081242300A787B3
0007240300912223
001126230007A483
00C1208300946C63
0041248300812403
0000806701010113
0004051300042783
000780E70047A783
0004222300050463
FCDFF06F00C40413
000037B7FF010113
000034B700912223
0011262300812423
0121202393478413
9704849393478793
0005091300941C63
0294146300078413
0440006F00000413
0007086300442703
0007270300042703
00C4041302A70863
00442783FD1FF06F
00C4041300079663
00042783FCDFF06F
0007A58300090513
FE0514E3D19FF0EF
00C1208300040513
0041248300812403
0101011300012903
0080079300008067
0000006F3007B7F3
00112623FF010113
FE010113FEDFF0EF
00112E2300912A23
0005049300812C23
7A0000EF00B12623
0005041300C12583
FCDFF0EF00048513
0181240300040513
0141248301C12083
1E10006F02010113
000037B700003537
AB87879398850613
0000059340C78633
CA1FF06F98850513
00200513FF010113
E71FF0EF00112623
000035B700003637
8786061300003537
8D8505138B858593
00300513F2CFF0EF
0A1000EFE4DFF0EF
000037B7FB5FE0EF
00C7C703A1C78793
00E78623FFE77713
0101011300C12083
F601011300008067
000047B708812C23
0931262300003437
A8C409938C078793
0101079300F9A223
0000059307000613
08112E2300078513
0921282308912A23
C01FF0EF09412423
00A9A42300100A13
01410EA300000513
00100513DCDFF0EF
10100793DC5FF0EF
670000EF00F11E23
00003937000037B7
000016B790078793
A1C90493000035B7
0000071300F12223
0141202300000793
0000081300000893
400006136E868693
A1C90513AC058593
718000EF0299A023
A8C4041300D4C783
00E486A3FFB7F713
00079A6301B7F793
000796630184A783
308000EFA1C90513
90878793000037B7
0000353700F12223
000026B700100793
9AC50493000035B7
00F0089300F12023
0000079300000813
4906869300000713
EC05859320000613
6A8000EF9AC50513
0094262300D4C783
FFB7F79300800513
000037B700F486A3
00F42C23AA478793
3005357300F42E23
9B1FE0EF00857513
0005278300452703
00E7A22300F72023
0005222300052023
00D5478300008067
0007986301F7F793
0015351301852503
0000051300008067
FF01011300008067
0000343700812423
000427839A440413
0207886300112623
0004278393DFF0EF
00C1208300812403
0000373700A78533
00000593A8A72E23
0101011300078513
00C120832050006F
0101011300812403
FF01011300008067
0011262300812423
3004347300800413
A807AE23000037B7
00A0079300950513
000037B702F55533
9AA7A22300847413
9AB7A023000037B7
30042473F6DFF0EF
0081240300C12083
0000806701010113
00812423FF010113
0011262300912223
0080041300050493
EFDFF0EF30043473
0084741300D4C783
00F486A3FFD7F793
00C1208330042473
0004A42300812403
0101011300412483
0085F79300008067
0000373700078C63
00071663A8C72703
861FE06F00058513
000080673007A7F3
00078A6300857793
A8C7270300003737
841FE06F00071463
000080673007A7F3
3005357300800513
FD5FF06F00857513
3007B7F300800793
A947268300003737
FFF7071300F6C703
0087F79300E687A3
000080673007A7F3
00F5146300052783
0007851300000793
FE01011300008067
0000343700812C23
0005049300912A23
02450513A8C40513
FCDFF0EF00112E23
00051463A8C40413
0084278300C42503
00D7C70302049A63
0207146301F77713
07F0071300E7D683
02F4202300D77E63
0181240301C12083
0201011301412483
00F5086300008067
E09FF0EF00A12623
02A4202300C12503
FF010113FD9FF06F
0011262300812423
3004347300800413
A947A703000037B7
0084741300000513
0017879300F74783
F51FF0EF00F707A3
0081240330042473
0101011300C12083
FF010113EF1FF06F
0011262300812423
3004347300800413
A8C7079300003737
000036B70247A783
00847413AB068693
06D78063A8C70713
0287258304078E63
00E7880300E50603
0047A70305065063
00E5222300F52023
00A7A22300A72023
0407E79300D54783
0000051300F506A3
30042473ECDFF0EF
0081240300C12083
0000806701010113
0007A78300B78663
02872783FA079AE3
00F5222300D52023
00A7A02302872783
FB5FF06F02A72423
FF010113FF052783
0121202300812423
0091222300112623
FE85091300050413
0080049302078663
000905133004B4F3
FF544783C99FF0EF
FFD7F7930084F493
3004A4F3FEF40AA3
FF544783FE042823
FEB7F79300090513
C89FF0EFFEF40AA3
0081240302050063
0041248300C12083
0001290300090513
ED9FF06F01010113
0081240300C12083
0001290300412483
0000806701010113
00812423FF010113
0011262300912223
0080049300050413
00D547833004B4F3
0407F7930084F493
C05FF0EF00078463
A8C7069300003737
0286A6030246A783
AB068693000036B7
06D78463A8C70713
00E4058306078263
04A5D66300E78503
00F420230047A683
0086A02300D42223
00D447830087A223
0407E79300872503
00F406A340850533
D69FF0EF00153513
00C120833004A4F3
0041248300812403
0000806701010113
0007A78300C78663
00C42223FA0794E3
00D4202302872783
028724230087A023
000037B7FADFF06F
000037B79A47A703
06070463A8C78793
07F006930087A703
04C6EC6300E75603
00E70603000036B7
04D644639A06A683
9AC6061300003637
0187268302C70E63
0107A68302069A63
FF01011302D54063
0011262300070513
00C12083ED9FF0EF
B39FF06F01010113
00D7A82340A686B3
0007A82300008067
FF01011300008067
0091222300812423
0005049300112623
3004347300800413
0084741300D54783
00078A630407F793
00D4C783AB9FF0EF
00F486A3FBF7F793
A947A503000037B7
0015351340950533
30042473C5DFF0EF
0081240300C12083
0101011300412483
000037B700008067
02478713A8C78793
02E7A42302E7A223
0000051300000593
000037B7AF5FF06F
00008067A947A503
01F7F79300D54783
0185250300079863
0000806700153513
0000806700000513
00812423FF010113
0091222300112623
3004347300800413
0084741300D54783
00071E630047F713
00C1208330042473
0041248300812403
0000806701010113
00F506A3FFB7F793
F95FF0EF00050493
0004851300050663
00040593C65FF0EF
00C1208300812403
0000353700412483
01010113AB850513
00400793AEDFF06F
00F506A300E50623
000507A300D50723
00052E2300052C23
0605202304052E23
FE01011300008067
00812C2302012303
0061202300112E23
B98FF0EF00050413
A947A783000037B7
0687A78301C12083
0181240306F42423
0000806702010113
FF01011306052783
0011262300812423
0007846300050413
00040513000780E7
02050463EE1FF0EF
E41FF0EF00040513
00C1208300D44783
00F406A30087E793
0101011300812403
00D4478300008067
000786630027F793
9DDFF0EF00040513
FC0786E301842783
2F4000EF01840513
FD010113FC1FF06F
03212023000037B7
0281242300003937
0211262302912223
01412C2301312E23
9707849397078413
03246E6397090913
A2DFF0EF00048413
00A00993FFF00493
0724646300002A37
02C1208302812403
0201290302412483
01812A0301C12983
AB9FF06F03010113
00F1222302C42783
00F1202302042783
01C4288301442783
0104270301842803
0084260300C42683
0004250300442583
00042783EB5FF0EF
030404130487AE23
02442603F85FF06F
0004250300960863
DEDFF0EF00061863
F81FF06F03040413
0336563300960613
01850513BD0A0593
12C000EF00160613
FD010113FE1FF06F
0211262302812423
0080059300050413
0085F5933005B5F3
E85FF0EF00B12623
A8C78793000037B7
00C125830087A703
0007A78302871263
0005851300079E63
02C1208395CFE0EF
0301011302812403
01C1051300008067
FE9FF06F8CDFF0EF
9A87A783000037B7
918FF06F00079463
0000806700000513
0205026300052783
9287270300003737
00078A6300E50C63
008526830087A703
00E7A42300D70733
00F7202300452703
0005202300E7A223
0000806700052223
FF010113000037B7
0081242392478793
001126230007A403
0000041300F41463
02040C63F89FF0EF
40A7853300842783
0000051300055463
A9C7A783000037B7
00A7D46300078663
00C1208300078513
0101011300812403
8000053700008067
FD5FF06FFFF54513
00812C23FE010113
00112E2300912A23
00C1262300050413
0080049300B52623
F1DFF0EF3004B4F3
0084F49300C12603
0010061300C04463
9247A703000037B7
00C4242300A60633
00F7066392478793
020710630047A583
00F420230047A703
0047A70300E42223
0087A22300872023
0087260302C0006F
04C6D86300842683
00D7242340D606B3
00E4202300472683
0086A02300D42223
0007A70300872223
00E4186300F70A63
00000593EF1FF0EF
3004A4F3FB1FE0EF
0181240301C12083
0201011301412483
40C686B300008067
F8B702E300D42423
F79FF06F00072703
00812423FF010113
0080041300112623
0005278330043473
0207806300847413
00000513E59FF0EF
00C1208330042473
0101011300812403
FEA0051300008067
FF010113FE9FF06F
0081242300112623
3007B47300800793
00847793E61FF0EF
00C120833007A7F3
0101011300812403
FE01011300008067
00912A2300812C23
0005049300112E23
0080041300B12623
E25FF0EF30043473
0084741300100793
00C1258300A7DA63
0004851300A4D663
30042473ED1FE0EF
0181240301C12083
0201011301412483
FE01011300008067
00912A2300812C23
0121282300112E23
0141242301312623
0005049301512223
999FF0EF00800413
000039B730043473
0000393700003A37
008474139A99A423
924A0A139A898993
00800A9399090913
0009A783000A2483
0049250300092683
00048A6301448C63
06E7D0630084A703
00E4A42340F70733
41F7D71300D786B3
00F6B7B300A70733
00D9202300E787B3
0009A02300F92223
00000593D51FF0EF
30042473E11FE0EF
0181240301C12083
0101290301412483
00812A0300C12983
0201011300412A83
00D706B300008067
00A585B341F75593
00B6063300E6B633
0004A42340E787B3
00D9202300048513
00F9A02300C92223
30042473CB1FF0EF
0004851300C4A783
300AB473000780E7
F3DFF06F00847413
00812423FF010113
0080041300112623
E49FF0EF300437F3
0010051300A04463
E69FF0EF00100593
FE5FF06FD7DFE0EF
00812423FF010113
0000343700912223
00112623000034B7
9704849397040413
00C1208300946E63
0041248300812403
0101011300000513
0144079300008067
00F42A2300040513
9DCFE0EF00F42C23
FCDFF06F01C40413
0000000000008067
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
00000000000010D4
0000000000001264
0000000000001264
0000000000001264
0000000000000FDC
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000000000001264
0000287800001264
0000000000000F20
00000F5000002878
0000288400000000
00000000000011DC
000014200000287C
000028780000292C
00000000000024C0
0303030302020100
0404040404040404
0505050505050505
0505050505050505
0606060606060606
0606060606060606
0606060606060606
0606060606060606
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
666C6F7672657773
0000737978656E5F
6F57206F6C6C6548
0A73252021646C72
7472617500000000
5F73797300000030
0000006B636F6C63
0000152C00001500
000000000000154C
0000293400000000
0000297000002964
0000297000002970
762D72796870657A
37312D302E312E32
3130316635672D33
0038303432373435
746F6F42202A2A2A
6870655A20676E69
756220534F207279
2520732520646C69
00000A2A2A2A2073
000000006E69616D
00000000656C6469
0001C20080002000
000007D000000000
000029240000140C
02FAF08000002924
0000274CFFFFFFF5
0000000000000000
0000000000002728
0000274000000000
0000291000002890
000000000000271C
0000273400000000
0000000000000000
0000297000002970
0000000000000000
000000000000000F
