0000000000000067
