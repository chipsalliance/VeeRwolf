0102829300000297
5080006F30529073
00112023FB010113
0041242300312223
0061282300512623
01C12C2300712A23
03E1202301D12E23
02A1242303F12223
02C1282302B12623
02E12C2302D12A23
0501202302F12E23
341022F305112223
300022F304512423
1F0000EF04512623
02051E6300000313
800003B7342022F3
0072F2B3FFF38393
00628A6300B00313
0000009700010513
3B00006F13408093
0042829304812283
0900006F04512423
0000239700010293
0043A10345838393
00512023FF010113
001E0E130003AE03
0003086301C3A023
03C0809300000097
342025733F80006F
FFF28293800002B7
158000EF00557533
E702829300002297
00A282B300351513
0042A3030002A503
00002317000300E7
000323833F830313
00732023FFF38393
0002811300012283
02032E0300832383
00002297087E0863
0082A3033D028293
0293282302832623
03332C2303232A23
0553202303432E23
0573242305632223
0593282305832623
05B32C2305A32A23
0000239702232423
0003AE0324038393
0202A30307C32623
028321030062A423
0303248302C32403
0383298303432903
04032A8303C32A03
04832B8304432B03
05032C8304C32C03
05832D8305432D03
3412907304812283
3002907304C12283
0041218300012083
00C1228300812203
0141238301012303
01C12E8301812E03
02412F8302012F03
02C1258302812503
0341268303012603
03C1278303812703
0441288304012803
3020007305010113
0000229700000073
0082A3032E028293
0085751306C32383
00038513300522F3
0010031300008067
3442B37300A312B3
342022F300008067
0062F2B380000337
0002846300000513
0000806700150513
0200079302060063
00F04C6340C787B3
00000713FE060513
0007059300A5D533
00C5D73300008067
00F595B300C55533
FE9FF06F00B56533
00002537000025B7
FE850513FD858593
FF0101132DD0006F
0081242300112623
02F5046300600793
020504635D8010EF
040516635D0010EF
2AC58593000025B7
2C05051300002537
2E1000EF2A5000EF
5BC010EFFFDFF06F
00002437FC051CE3
0084258350C40413
2E05051300002537
0084250327D000EF
FD1FF06F7DC010EF
2A858593000025B7
FB010113FB9FF06F
0491222304812423
0060079304112623
0005841300050493
000027370EA7E063
FFC7071300251793
0007A78300E787B3
0000253700078067
221000EF12C50513
04442783504010EF
00C4280301042883
0404278302F12823
0004268300442703
03C4278302F12623
0005059304842603
0384278302F12423
1B05051300002537
0344278302F12223
0304278302F12023
02C4278300F12E23
0284278300F12C23
0244278300F12A23
0204278300F12823
01C4278300F12623
0184278300F12423
0144278300F12223
0084278300F12023
0004059318D000EF
EA9FF0EF00048513
1545051300002537
00002537F55FF06F
F49FF06F17050513
0004859300002537
159000EF18C50513
FF010113F39FF06F
0011262300812423
3420267300050413
0016561300161613
02C7E86300500793
0026179300002737
00F707B301870713
000025370007A583
111000EF03850513
0000051300040593
000025B7EA5FF0EF
FE1FF06F03058593
00112623FF010113
00002537342025F3
0015D59300159593
0D9000EF30850513
05458593000025B7
E69FF0EF00400513
41078793000027B7
00070C630007A703
0007A0230007A303
4147A503000027B7
0000806700030067
00112623FF010113
101000EF455000EF
000021174B9000EF
000012B762C10113
0051013380028293
21C0006FFD9FF0EF
01312E23FD010113
0301268300068993
0321202302812423
0006091300058413
0040061300088593
0211262302912223
00E1262300050493
0101222300F12423
00812783578010EF
00B405B3FB090593
0604A0230404AE23
02F5A823FF05F593
00C12703000027B7
8807879300412803
000007B704F5A623
0281240302C12083
0335A42352C78793
0305AA2302E5A623
02B4A42304F5A423
0241248302012903
0301011301C12983
00C0079300008067
00C5278302F58733
00B5070300E787B3
0007A78300B75463
02E6473302000713
0027171301F67513
00F6A02300E787B3
FE01011300008067
00112E2300C10693
00C12703FBDFF0EF
00A7953300100793
01C1208300072783
00F7202300A7E7B3
0000806702010113
0085580300452783
00812423FF010113
0005041302F80833
00A4488300052503
00112623FFF00713
00E405A300912223
00C0031300000593
01F00E1301050533
0315C26302000E93
0084578300000493
00C1208306F4C463
0041248300812403
0000806701010113
00C4260302F85733
00D606B3026586B3
00C6A22300468613
00EE4E6300C6A423
0027D79300B405A3
FFC7F79300378793
FA9FF06F00158593
03D7473301F70713
0027171300A6A023
FD9FF06F00E50533
0004861300442783
02F4873300000593
0004051300042783
00E787B300148493
0047069300C42703
0087268300D7A023
0087268300D7A223
00F7242300F6A023
F51FF06FED5FF0EF
00050793FF010113
0006059300058513
0011262300068613
120010EF000780E7
0000051339C010EF
FF01011300008067
0005041300812423
0011262304500513
0005849300912223
00048593000400E7
000400E705200513
0081240300040313
0004859300C12083
0520051300412483
0003006701010113
001787930005A783
000027B700F5A023
000300673AC7A303
04812423FB010113
03412C2303312E23
0361282303512A23
0491222304112623
0371262305212023
0391222303812423
01B12E2303A12023
00058A9300050A13
00068B1300060993
00E0546300100413
0010079300070413
00FB146302000C13
3B9AD4B703000C13
00A00C9300100913
9FF4849300000713
00A00D1300200D93
0007146300148B93
0379D5330934F263
00190913000A8593
000A00E703050513
FFFC8C9300100713
0379F9B300100793
FCFC96E303A4D4B3
03098513000A8593
00300793000A00E7
06FB0A6341240433
0481240304C12083
0401290304412483
03812A0303C12983
03012B0303412A83
02812C0302C12B83
02012D0302412C83
0501011301C12D83
F9944CE300008067
000A8593F96DEAE3
00E12623000C0513
00190913000A00E7
F79FF06F00C12703
02000513000A8593
FFF40413000A00E7
F8DFF06FFE8048E3
3AA7A623000027B7
FB01011300008067
0491222304812423
03312E2305212023
03512A2303412C23
03A1202303912223
0411262301B12E23
0371262303612823
0005041303812423
00060A9300058493
00000A1300068D13
00000993FFF00913
80000DB700000C93
04051063000AC503
0481240304C12083
0401290304412483
03812A0303C12983
03012B0303412A83
02812C0302C12B83
02012D0302412C83
0501011301C12D83
000C9E6300008067
36D50A6302500693
000400E700048593
FA5FF06F001A8A93
10D50E6306400693
0390069306A6E263
0310069302A6EA63
02D006930ED57463
0300079334D50A63
025007130CF50063
0004859302E51263
000400E702500513
0580069315C0006F
063007131AD50E63
000485932EE50E63
000400E702500513
000AC50300048593
07000693FD5FF06F
02A6E06316D50A63
0AD5026306900693
08D50A6306C00693
F6D506E306800693
07500693FC5FF06F
02A6EE6310D50663
FAE518E307300713
004D0B13000D2C03
000BC503000C0B93
0030079326051863
418B8BB300F99863
2770466341790BB3
0C80006F000B0D13
12D5046307800693
FA9FF06F07A00693
2809886300095E63
F00992E3FD050913
EFDFF06F00200993
00A00693FE0948E3
FD09091302D90933
FE1FF06F01250933
EDDFF06F001A0A13
000D2603040A1263
02065063004D0D13
02D0051300048593
000400E700C12023
FFF9091300012603
0009071340C00633
0004859300098693
C95FF0EF00040513
0010071303C0006F
007D0793FAEA0EE3
00072603FF87F713
00870D1300472683
00C7373301B60733
FA0700E300D70733
0004051300048593
00000C93BF5FF0EF
000A1863E59FF06F
004D0D13000D2603
00100713F9DFF06F
007D0793FEEA08E3
00870D13FF87F713
0047270300072603
800007B7FC0710E3
F6C7F8E3FFF7C793
00048593FB1FF06F
000400E703000513
0780051300048593
00800913000400E7
0010069300100993
000D27830B46C263
004D0D1300012423
01000C1300F12223
0001202300000B93
0041250301000893
FFF88B1300812583
01112623002B1613
00F57513E50FF0EF
0001278308051863
0007986303000693
0010079300C12883
00A6853308F89663
0004859301851513
000400E741855513
040B1863001B8B93
00000C9300300693
00191713D6D998E3
F17054E341770BB3
0200051300048593
FFFB8B93000400E7
007D0793FEDFF06F
0006A783FF87F693
00F1222300868D13
00F124230046A783
01912023F55FF06F
F59FF06F000B0893
0570069300900793
03000693F8A7E2E3
FFFC0793F7DFF06F
01894C6300F12623
00F99C6300100793
0300051300048593
00C12C03000400E7
00200793FC1FF06F
00048593FEF99AE3
FE5FF06F02000513
001B8B9300048593
D81FF06F000400E7
0200051300048593
FFFB8B93000400E7
000D2503D85FF06F
004D0B1300048593
D75FF06F000400E7
FFF0091300000A13
00100C9300000993
00300993C89FF06F
00100993C81FF06F
FE010113C79FF06F
0000053700050613
7C05051300058693
00112E2300C10593
BA1FF0EF00012623
0201011301C12083
FC01011300008067
0241059302B12223
02C1242300112E23
02E1282302D12623
03012C2302F12A23
00B1262303112E23
01C12083FA5FF0EF
0000806704010113
0080079300008067
105000733007A7F3
0010079300008067
3045257300A79533
0010079300008067
3045357300A79533
0080079300008067
304050733007B7F3
0000806734405073
00812423FF010113
0000243700912223
00A0079300112623
4184041300050493
0004250300F51C63
0045278300D00593
000780E70047A783
0FF4F59300042503
0047A78300452783
00C12083000780E7
0004851300812403
0101011300412483
FF01011300008067
0000143700812423
00112623E2040513
E2040513188000EF
00C1208300812403
A75FF06F01010113
FF01011300002537
0011262333050513
000027B7200000EF
FB9FF0EF40A7AC23
0000051300C12083
0000806701010113
00700513FF010113
F11FF0EF00112623
0186A783800016B7
090707130003D737
0070051300E787B3
EE1FF0EF00F6AC23
0010051300C12083
6A50006F01010113
00700513FF010113
ED1FF0EF00112623
0186A783800016B7
090707130003D737
0070051300E787B3
EA1FF0EF00F6AC23
0000051300C12083
0000806701010113
0000051300008067
0005478300008067
00E794630005C703
40E7853300079663
0015051300008067
FE1FF06F00158593
000507930FF5F693
040718630037F713
008597130FF5F593
0105971300B765B3
00C7833300B765B3
0030081300078713
03186E6340E308B3
0027159300265713
FFC0059300B787B3
00C7073302B70733
02E7946300E78733
FE060EE300008067
FED78FA300178793
F9DFF06FFFF60613
FEB72E2300470713
00178793FB9FF06F
FD1FF06FFED78FA3
00008067FFF00513
3AA7A823000027B7
800017B700008067
0000806700B78423
0087C783800017B7
00F5802300000513
0000051300008067
0025171300008067
00150513000027B7
0025151335878793
00E78733FF010113
0081242300A787B3
0007240300912223
001126230007A483
00C1208300946C63
0041248300812403
0000806701010113
0004051300042783
000780E70047A783
0004222300050463
FCDFF06F00C40413
000027B7FF010113
000024B700912223
0011262300812423
012120233C478413
3F4484933C478793
0005091300941C63
0294146300078413
0440006F00000413
0007086300442703
0007270300042703
00C4041302A70863
00442783FD1FF06F
00C4041300079663
00042783FCDFF06F
0007A58300090513
FE0514E3E35FF0EF
00C1208300040513
0041248300812403
0101011300012903
0000253700008067
40850613000027B7
40C7863353878793
4085051300000593
FF010113E19FF06F
0011262300200513
00002537ECDFF0EF
C09FF0EF36C50513
EB9FF0EF00300513
90CFF0EF061000EF
49C78793000027B7
FFE7771300C7C703
00C1208300E78623
0000806701010113
08812C23F6010113
00002437000037B7
3407879309312623
00F9A22350C40993
0700061301010793
0007851300000593
08912A2308112E23
D8DFF0EF09212823
00A9A42300100713
00E10EA300000513
00100513E3DFF0EF
10100793E35FF0EF
638000EF00F11E23
39C78793000027B7
00F1222300002937
00100793000016B7
49C90493000025B7
0000071300F12023
0000089300000793
17C6869300000813
5405859340000613
0299A02349C90513
00D4C7836D8000EF
FFB7F71350C40413
01B7F79300E486A3
0184A78300079A63
49C9051300079663
000027B72DC000EF
00F122233A478793
0010079300002537
000035B7000026B7
00F1202342C50493
0000081300F00893
0000071300000793
20000613EDC68693
42C5051394058593
00D4C783668000EF
0080051300942623
00F486A3FFB7F793
52478793000027B7
00F42E2300F42C23
0085751330053573
00452703F11FE0EF
00F7202300052783
0005202300E7A223
0000806700052223
01F7F79300D54783
0185250300079863
0000806700153513
0000806700000513
00112623FF010113
000027B7C05FF0EF
00C120834207A783
00A7853300002737
0000059350A72E23
0101011300078513
FF0101131E10006F
0011262300812423
3004347300800413
5007AE23000027B7
00A0079300950513
000027B702F54533
42A7A02300847413
40B7AE23000027B7
30042473F91FF0EF
0081240300C12083
0000806701010113
00812423FF010113
0011262300912223
0080041300050493
F21FF0EF30043473
0084741300D4C783
00F486A3FFD7F793
00C1208330042473
0004A42300812403
0101011300412483
000027B700008067
0007966350C7A783
DEDFE06F00058513
3005A5F30085F593
0000273700008067
0007146350C72703
00857793DD1FE06F
000080673007A7F3
3005357300800513
FD9FF06F00857513
3007B7F300800793
5147268300002737
FFF7071300F6C703
0087F79300E687A3
000080673007A7F3
00F5146300052783
0007851300000793
FE01011300008067
0000243700812C23
0005049300912A23
0245051350C40513
FCDFF0EF00112E23
0005146350C40413
0084278300C42503
00D7C70302049A63
0207146301F77713
07F0071300E7D683
02F4202300D77E63
0181240301C12083
0201011301412483
00F5086300008067
E35FF0EF00A12623
02A4202300C12503
FF010113FD9FF06F
0011262300812423
3004347300800413
5147A703000027B7
0084741300100513
0017879300F74783
F51FF0EF00F707A3
0081240330042473
0101011300C12083
FF010113EF1FF06F
0011262300812423
3004347300800413
50C7079300002737
000026B70247A783
0084741353068693
06D7806350C70713
0287258304078E63
00E7880300E50603
0047A70305065063
00E5222300F52023
00A7A22300A72023
0407E79300D54783
0000051300F506A3
30042473ECDFF0EF
0081240300C12083
0000806701010113
0007A78300B78663
02872783FA079AE3
00F5222300D52023
00A7A02302872783
FB5FF06F02A72423
FF010113FF052783
0121202300812423
0091222300112623
FE85091300050413
0080049302078663
000905133004B4F3
FF544783CC5FF0EF
FFD7F7930084F493
3004A4F3FEF40AA3
FF544783FE042823
FEB7F79300090513
CB5FF0EFFEF40AA3
0081240302050063
0041248300C12083
0001290300090513
ED9FF06F01010113
0081240300C12083
0001290300412483
0000806701010113
00812423FF010113
0011262300912223
0080049300050413
C41FF0EF3004B4F3
50C7079300002737
000026B70247A783
0084F49353068693
06D7866350C70713
0287258306078463
00E7850300E40603
0047A68304A65663
00D4222300F42023
0087A2230086A023
0087250300D44783
408505330407E793
0015351300F406A3
3004A4F3D75FF0EF
0081240300C12083
0101011300412483
00B7866300008067
FA0794E30007A783
00D4202302872783
0287278300F42223
028724230087A023
000027B7FA9FF06F
060786634207A783
50C78793000027B7
07F006930087A703
04C6EA6300E75603
00E70603000026B7
04D6426341C6A683
3C06A683000026B7
0187268302D70C63
0107A68302069863
FF01011302D54063
0011262300070513
00C12083EE1FF0EF
B6DFF06F01010113
00D7A82340A686B3
FF01011300008067
0091222300812423
0005049300112623
3004347300800413
0084741300D54783
00078A630407F793
00D4C783AF5FF0EF
00F486A3FBF7F793
5147A503000027B7
0015351340950533
30042473C6DFF0EF
0081240300C12083
0101011300412483
000027B700008067
0247871350C78793
02E7A42302E7A223
0000051300000593
000027B7B0DFF06F
000080675147A503
01F7F79300D54783
0185250300079863
0000806700153513
0000806700000513
50C7A503000027B7
0000806700A03533
5147A783000027B7
0015751300C7C503
FF01011300008067
0011262300812423
0080041300912223
00D5478330043473
0047F71300847413
3004247300071E63
0081240300C12083
0101011300412483
FFB7F79300008067
0005049300F506A3
00050663F71FF0EF
C51FF0EF00048513
0081240300040593
0041248300C12083
5385051300002537
AE1FF06F01010113
02012303FE010113
00112E2300812C23
0005041300612023
000027B7BC9FE0EF
01C120835147A783
06F424230687A783
0201011301812403
0605278300008067
00812423FF010113
0005041300112623
000780E700078463
EE5FF0EF00040513
0004051302050463
00D44783E45FF0EF
0087E79300C12083
0081240300F406A3
0000806701010113
0027F79300D44783
0004051300078663
018427839F9FF0EF
01840513FC0786E3
FC1FF06F2FC000EF
000027B7FD010113
0000293703212023
0291222302812423
01312E2302112623
3F47841301412C23
3F4909133F478493
0004841303246E63
FFF00493A41FF0EF
00001A3700A00993
0281240307246463
0241248302C12083
01C1298302012903
0301011301812A03
02C42783ACDFF06F
0204278300F12223
0144278300F12023
0184280301C42883
00C4268301042703
0044258300842603
EB5FF0EF00042503
0487AE2300042783
F85FF06F03040413
0096086302442603
0006186300042503
03040413E15FF0EF
00960613F81FF06F
628A059303364633
0016061301850513
FE1FF06F134000EF
00C506A300D50623
000507A300B50723
00052E2300052C23
FD01011300008067
0080059302112623
0085F5933005B5F3
E71FF0EF00B12623
01C1051300C12583
02C12083905FF0EF
0000806703010113
4247A783000027B7
C20FF06F00079463
0000806700000513
0205026300052783
3B87270300002737
00078A6300E50C63
008526830087A703
00E7A42300D70733
00F7202300452703
0005202300E7A223
0000806700052223
4287C783000027B7
00112623FF010113
0091222300812423
00079663FFF00513
FFF5451380000537
3B478793000027B7
02F404630007A403
0084248302040263
40A484B3F69FF0EF
0004C86300000513
F55FF0EF00842403
000027B740A40533
0007866351C7A783
0007851300A7D463
0081240300C12083
0101011300412483
FE01011300008067
00912A2300812C23
0005041300112E23
00B5262300C12623
3004B4F300800493
00C12603F01FF0EF
00C044630084F493
000027B700100613
00A606333B47A703
3B47879300C42423
0047A58300F70663
0047A70302071063
00E4222300F42023
008720230047A703
02C0006F0087A223
0084268300872603
40D606B304C6D863
0047268300D72423
00D4222300E42023
008722230086A023
00F70A630007A703
ED5FF0EF00E41863
A9CFF0EF00000593
01C120833004A4F3
0141248301812403
0000806702010113
00D4242340C686B3
00072703F8B702E3
FF010113F79FF06F
0011262300812423
3004347300800413
0084741300052783
E3DFF0EF02078063
3004247300000513
0081240300C12083
0000806701010113
FE9FF06FFEA00513
00112623FF010113
0080079300812423
E45FF0EF3007B473
3007A7F300847793
0081240300C12083
0000806701010113
00812C23FE010113
00112E2300912A23
00B1262300050493
3004347300800413
00847413E09FF0EF
00A4DA6300C12583
00A7D66300100793
9BCFF0EF00048513
01C1208330042473
0141248301812403
0000806702010113
00812C23FE010113
00112E2300912A23
0131262301212823
0151222301412423
0080041300050493
3004347399DFF0EF
00002A37000029B7
4299A22300002937
4249899300847413
408909133B4A0A13
000A248300800A93
000926830009A783
01448C6300492503
0084A70300048A63
40F7073306E7D063
00D786B300E4A423
00A7073341F7D713
00E787B300F6B7B3
00F9222300D92023
D35FF0EF0009A023
8FCFF0EF00000593
01C1208330042473
0141248301812403
00C1298301012903
00412A8300812A03
0000806702010113
41F7559300D706B3
00E6B63300A585B3
40E787B300B60633
000485130004A423
00C9222300D92023
C95FF0EF00F9A023
00C4A78330042473
000780E700048513
00847413300AB473
FF010113F3DFF06F
0011262300812423
300437F300800413
00A04463E49FF0EF
0010059300100513
ED9FE0EFE69FF0EF
FF010113FE5FF06F
0091222300812423
000024B700002437
3F44041300112623
00946E633F448493
0081240300C12083
0000051300412483
0000806701010113
0004051301440793
00F42C2300F42A23
01C40413EF0FE0EF
00008067FCDFF06F
000004A800000000
000004A800000000
000004A800000000
000004A800000000
000004A800000000
000004A800000000
000004A800000000
00000EE000000000
00000EB000002050
0000233800000000
0000000000000F20
0000104C00002330
0000205000000000
0000000000001F0C
666C6F7672657773
0000737978656E5F
6F57206F6C6C6548
0A73252021646C72
0000038000000000
0000043800000438
0000038000000374
0000042C00000420
000020C4000020A4
000020F4000020E0
0000211800002100
006E776F6E6B6E75
6F69747065637845
206573756163206E
0A29642528207325
DEADBAAD00000000
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
74736E49DEADBAAD
206E6F6974637572
2073736572646461
6E67696C6173696D
74736E4900006465
206E6F6974637572
6620737365636341
00000000746C7561
206C6167656C6C49
7463757274736E69
61657242006E6F69
0000746E696F706B
6464612064616F4C
73696D2073736572
0064656E67696C61
6363612064616F4C
6C75616620737365
2A2A2A2A00000074
206C656E72654B20
697461636F6C6C41
756C696146206E6F
2A2A2A2A20216572
2A2A2A2A0000000A
6C656E72654B202A
2A202153504F4F20
0000000A2A2A2A2A
654B202A2A2A2A2A
6E6150206C656E72
2A2A2A2A20216369
2A2A2A2A00000A2A
6E776F6E6B6E5520
45206C6174614620
21642520726F7272
00000A2A2A2A2A20
20746E6572727543
4920646165726874
460A7025203D2044
20676E69746C7561
7463757274736E69
72646461206E6F69
7830203D20737365
3A617220200A7825
6720207825783020
2078257830203A70
257830203A707420
30203A3074202078
317420200A782578
202078257830203A
78257830203A3274
7830203A33742020
203A347420207825
7420200A78257830
2078257830203A35
257830203A367420
30203A3061202078
3A31612020782578
20200A7825783020
78257830203A3261
7830203A33612020
203A346120207825
3561202078257830
200A78257830203A
257830203A366120
30203A3761202078
000000000A782578
6573736500525349
6874206C6169746E
0000000064616572
6166206C61746146
25206E6920746C75
6E6E697053202173
000A2E2E2E676E69
6166206C61746146
74206E6920746C75
7025206461657268
6974726F62412021
000000000A2E676E
73756F6972757053
75727265746E6920
6365746564207470
5152492021646574
0000000A6425203A
0000003074726175
636F6C635F737973
000010380000006B
000000000000102C
0000000000000000
000023E8000023C4
000023F4000023F4
2A2A2A2A000023F4
6E69746F6F42202A
72796870655A2067
6870657A20534F20
34312E31762D7279
2A2A2A2A2A20302E
6E69616D0000000A
656C646900000000
0000076C00000000
000023B400001018
FFFFFFF5000023B4
00001FCC0000242C
0000000000000000
0000234400001FC0
00001FA800000000
0000000000000000
0000000000001FB4
000023F400000000
00000000000023F4
0000000F00000000
