0102829300000297
47D0006F30529073
00112023FB010113
0041242300312223
0061282300512623
01C12C2300712A23
03E1202301D12E23
02A1242303F12223
02C1282302B12623
02E12C2302D12A23
0501202302F12E23
341022F305112223
300022F304512423
1F0000EF04512623
02051E6300000313
800003B7342022F3
0072F2B3FFF38393
00628A6300B00313
0000009700010513
3250006F13408093
0042829304812283
0900006F04512423
0000639700010293
0043A10345C38393
00512023FF010113
001E0E130003AE03
0003086301C3A023
03C0809300000097
3420257336D0006F
FFF28293800002B7
158000EF00557533
4382829300005297
00A282B300351513
0042A3030002A503
00006317000300E7
000323833FC30313
00732023FFF38393
0002811300012283
02032E0300832383
00006297087E0863
0082A3033D428293
0293282302832623
03332C2303232A23
0553202303432E23
0573242305632223
0593282305832623
05B32C2305A32A23
0000639702232423
0003AE03F1038393
0202A30307C32623
028321030062A423
0303248302C32403
0383298303432903
04032A8303C32A03
04832B8304432B03
05032C8304C32C03
05832D8305432D03
3412907304812283
3002907304C12283
0041218300012083
00C1228300812203
0141238301012303
01C12E8301812E03
02412F8302012F03
02C1258302812503
0341268303012603
03C1278303812703
0441288304012803
3020007305010113
0000629700000073
0082A3032E428293
0085751306C32383
00038513300522F3
0010031300008067
3442B37300A312B3
342022F300008067
0062F2B380000337
0002846300000513
0000806700150513
0200079302060063
00F04C6340C787B3
00000713FE060513
0007059300A5D533
00C5D73300008067
00F595B300C55533
FE9FF06F00B56533
0006081300058793
0005031300068893
0000573728069663
0EC5F6635A070713
0CD67863000106B7
00C6B6B30FF00693
00D658B300369693
0007470301170733
0200071300D706B3
00070C6340D70733
00D556B300E797B3
00F6E5B300E61833
0108551300E51333
0108161302A5F733
0103569301065613
0107171302A5D5B3
02B607B300D766B3
00F6FE6300058713
FFF58713010686B3
00F6F6630106E863
010686B3FFE58713
02A6F7B340F686B3
0103531301031313
0107979302A6D6B3
02D605B30067E333
00B37C6300068513
FFF6851300680333
00B3746301036663
01071713FFE68513
0000059300A76733
010008B70E40006F
F3166CE301000693
F31FF06F01800693
0010069300061663
000106B702C6D833
0FF006930CD87263
008008930106F463
00D70733011856B3
0200071300074683
40D70733011686B3
410787B30A071863
0108561300100593
0108D89301081893
02C7F73301035693
0107171302C7D7B3
02F8853300D766B3
00A6FE6300078713
FFF78713010686B3
00A6F6630106E863
010686B3FFE78713
02C6F7B340A686B3
0103531301031313
0107979302C6D6B3
02D888B30067E333
01137C6300068513
FFF6851300680333
0113746301036663
01071713FFE68513
0007051300A76733
010006B700008067
F4D862E301000893
F3DFF06F01800893
00D7D5B300E81833
00D556B300E51333
00E797B301085513
00F6E8B302A5F733
0107D79301081793
02A5D5B30108D613
00C7673301071713
0005861302B786B3
0107073300D77E63
01076863FFF58613
FFE5861300D77663
40D706B301070733
0108989302A6F733
02A6D6B30108D893
02D785B301071713
00068713011767B3
010787B300B7FE63
0107E863FFF68713
FFE6871300B7F663
40B787B3010787B3
00E5E5B301061593
18D5E663EB5FF06F
04E6F46300010737
00D837330FF00813
0000583700371713
00E6D5B35A080813
0005C803010585B3
00E8083302000593
02059663410585B3
EEF6ECE300100713
0015471300C53533
010005B7EEDFF06F
FCB6E0E301000713
FB9FF06F01800713
00B696B301065733
0106DE9300D766B3
03D778B30107D733
0105583300B797B3
0106979300F86333
010358130107D793
03D7573300B61633
0108E83301089893
00070E1302E78F33
00D8083301E87E63
00D86863FFF70E13
FFE70E1301E87663
41E8083300D80833
03D8583303D878B3
03078EB301089893
0107D79301031793
0008071300F8E7B3
00D787B301D7FE63
00D7E863FFF80713
FFE8071301D7F663
010E1E1300D787B3
00010EB741D787B3
FFFE881300EE6733
0107589301077333
0106561301067833
0308883303030E33
02C30333010E5693
006686B301030333
0106F46302C888B3
0106D61301D888B3
0317E663011608B3
000107B7CF179AE3
00F6F6B3FFF78793
00FE7E3301069693
01C686B300B51533
DAD57CE300000593
CC9FF06FFFF70713
0000071300000593
FE010113DA5FF06F
00812C2300112E23
0006041300912A23
0121282300058493
6AD030EF00050913
00A126232DD030EF
0010061300006537
8905051300190593
00C12703091010EF
0000663706074263
88C60613000066B7
000065378B468693
89C5051300090593
06040063069010EF
0487D6633E700793
90C58593000065B7
0004851300040613
01812403049010EF
0141248301C12083
0000653701012903
02010113A0C50513
000066370290106F
88860613000066B7
FA1FF06F90C68693
8B458593000065B7
000065B7FB9FF06F
0004851390C58593
FB1FF06F7F8010EF
02912A23FC010113
02112E2303412423
0321282302812C23
0351222303312623
01712E2303612023
01912A2301812C23
01B1262301A12823
0005049300500793
0EF50E6300150A13
6A078793000057B7
00E7873300251713
002A171300072903
0007A98300E787B3
00006D3700006DB7
01900A9306400B13
00006C3700006CB7
0000061300006BB7
00048513810D8593
FFF00593E95FF0EF
164020EF00090513
828D059300000613
E79FF0EF00048513
00098513FFF00593
429040EF148020EF
840C859303655433
0344043300048513
0014041301F47413
0004061303540433
00040513E45FF0EF
00098513479030EF
858C059334C020EF
0004851300000613
00090513E25FF0EF
3D9040EF334020EF
870B859303655433
0344043300048513
0014041301F47413
0004061303540433
00040513DF5FF0EF
F49FF06F429030EF
1189099300006937
1189091306498993
00005637F19FF06F
00005537000055B7
6B860613FC010113
6C8505136C058593
02812C2302112E23
0321282302912A23
0341242303312623
0361202303512223
65C010EF01712E23
0000059300001537
594020EF38850513
1185041300006537
038020EF11850513
030020EF01440513
028020EF02840513
020020EF03C40513
018020EF05040513
0000693706440513
008020EF00006437
5509091319040413
00300A9300000493
00400B13FFF00B93
0060099300000A37
00048713409A88B3
0000081300090593
7C0A069300000793
0004051330000613
0161202301712223
00040513679030EF
545030EF00148493
3009091307040413
03C12083FD3490E3
0341248303812403
02C1298303012903
02412A8302812A03
01C12B8302012B03
0000806704010113
00112623FF010113
0060079300812423
391030EF02F50463
389030EF02050463
000065B704051663
00006537B6858593
544010EFB7C50513
FFDFF06F5B0010EF
FC051CE3375030EF
5104041300006437
0000653700842583
51C010EFB9C50513
7CD030EF00842503
000065B7FD1FF06F
FB9FF06FB6458593
04812423FB010113
0411262304912223
0005049300600793
0EA7E06300058413
0025179300006737
00E787B38B870713
000780670007A783
9E85051300006537
2BD030EF4C0010EF
0104288304442783
02F1282300C42803
0044270304042783
02F1262300042683
0484260303C42783
02F1242300050593
0000653703842783
02F12223A6C50513
02F1202303442783
00F12E2303042783
00F12C2302C42783
00F12A2302842783
00F1282302442783
00F1262302042783
00F1242301C42783
00F1222301842783
00F1202301442783
42C010EF00842783
0004851300040593
00006537EA9FF0EF
F55FF06FA1050513
A2C5051300006537
00006537F49FF06F
A485051300048593
F39FF06F3F8010EF
00812423FF010113
0005041300112623
0016161334202673
0050079300165613
0000673702C7E863
8D47071300261793
0007A58300F707B3
8F45051300006537
000405933B0010EF
EA5FF0EF00000513
8EC58593000065B7
FF010113FE1FF06F
342025F300112623
0015959300006537
BC4505130015D593
000065B7378010EF
0040051391058593
000067B7E69FF0EF
0007A7030E878793
0007A30300070C63
000067B70007A023
000300670EC7A503
FF01011300008067
2A1010EF00112623
305010EF3C0010EF
0C81011300007117
80028293000012B7
FD9FF0EF00510133
FD0101134BD0006F
0291222302812423
01312E2303212023
01512A2301412C23
0171262301612823
0211262300078B13
0280079301812423
0005841300050493
00068A1300060993
00080A9300070B93
08F89A6300088913
6E478793000027B7
0301268308F69A63
0004851300090593
19D030EF00400613
00B405B3FB098593
0404AE23000027B7
FF05F5930604A023
04F5A62388078793
02C12083000017B7
CA07879302812403
0375A6230345A423
0355AA230365A823
02B4A42304F5A423
0241248302012903
01812A0301C12983
01012B0301412A83
00812C0300C12B83
0000806703010113
0440079301D88693
00006C37F6D7FAE3
00006537000065B7
01800693BECC0613
C9850513C0C58593
00006537200010EF
FE30069300090593
CB85051302700613
018005931E8010EF
218010EFBECC0513
00C00793F2DFF06F
00C5278302F58733
00B5070300E787B3
0007A78300B75463
02E6473302000713
0027171301F67513
00F6A02300E787B3
FE01011300008067
00112E2300C10693
00C12703FBDFF0EF
00A7953300100793
01C1208300072783
00F7202300A7E7B3
0000806702010113
0085580300452783
00812423FF010113
0005041302F80833
00A4488300052503
00112623FFF00713
00E405A300912223
00C0031300000593
01F00E1301050533
0315C26302000E93
0084578300000493
00C1208306F4C463
0041248300812403
0000806701010113
00C4260302F85733
00D606B3026586B3
00C6A22300468613
00EE4E6300C6A423
0027D79300B405A3
FFC7F79300378793
FA9FF06F00158593
03D7473301F70713
0027171300A6A023
FD9FF06F00E50533
0004861300442783
02F4873300000593
0004051300042783
00E787B300148493
0047069300C42703
0087268300D7A023
0087268300D7A223
00F7242300F6A023
F51FF06FED5FF0EF
00C5222300058663
0005278300008067
00F666330017F793
0000806700C52023
FE01011300052783
00912A2300812C23
0131262301212823
0005099300112E23
00F6202300058913
0010049300060413
0325926300042583
0181240301C12083
0101290300048513
00C1298301412483
0000806702010113
000905130049A783
00042783000780E7
0047A78300051E63
FC0782E300440413
00F4202300148493
0007A783FB1FF06F
FE5FF06FFFE7F793
FD01011300259793
01612823FF878793
0321202300F50B33
00478793000B2903
00F504B302912223
0049278302812423
01412C230004A403
40F40A3301712623
01312E2302112623
001A3B9301512A23
00442A8308F41C63
08F40C6301403A33
0020079300442983
FFCB250300B7DE63
0045258300040613
0015B593412585B3
000A8613ED1FF0EF
00040513000B8593
00090613EC1FF0EF
00040513000A0593
00098613EB1FF0EF
00090513000B8593
02C12083EA1FF0EF
02812403008B2023
01C129830124A023
0201290302412483
01412A8301812A03
00C12B8301012B03
0000806703010113
FFEAFA9300042A83
00042983F69FF06F
F69FF06FFFE9F993
0005A7030085A783
0027969300178793
00D7073300F5A423
0045A70300A72023
00F707B300100693
0005250300078023
0005A7030085A783
00051A63FFE57513
00F707B300279793
000080670007A503
0027961300178793
00C7073300F5A423
0045A70300A72023
00D7802300F707B3
FD010113FBDFF06F
40000BB701712623
0161282301312E23
01A1202301812423
0281242302112623
0321202302912223
01512A2301412C23
00050D1301912223
00060B1300058993
FFFB8B9300100C13
01798A330F3C5863
014D0A33002A1A13
000A2903FFCA2483
41990AB30044AC83
000C8413001ABA93
0004A40301991663
00042783FFE47413
040790630017F793
008A202300098593
DF5FF0EF000D0513
001989930004A783
00F4A023FFE7F793
000A248300042783
00F420230017E793
07990463012A2223
00042A030044A403
FFEA7A1300442703
000A2783000A0863
140784630017F793
0007278300070863
080788630017F793
0000061301691A63
00048513000A8593
00042783CD9FF0EF
00F42023FFE7F793
0017F7130004A783
FFF9899300070C63
0004A403F29FF06F
F99FF06FFFE47413
00F4A0230017E793
0281240302C12083
0201290302412483
01812A0301C12983
01012B0301412A83
00812C0300C12B83
00012D0300412C83
0000806703010113
FFE7F79300042783
000A07931080006F
000707930B990863
0016F6930007A683
0004A7030A069263
0009859300042683
FFE6F69300177713
00E4202300D76733
000D05130004A703
00E4A02300176713
001767130007A703
0029979300E7A023
FE87AE2300FD07B3
F5691EE3CB1FF0EF
02C1208302812403
01C1298302012903
01012B0301812A03
00812C0300C12B83
00012D0300412C83
00048513000A8593
0241248301412A83
0301011300000613
000A0793BB9FF06F
00070793F79900E3
01991463F4079CE3
00299B9300070A13
017D0BB3FFCB8B93
014BA223008BA023
000D051300198593
00042783C31FF0EF
00F42023FFE7F793
000BA403000A2783
00FA20230017E793
00442783EF990CE3
F11FF06F012BA023
0005086300052503
0045278300058C63
0000806700079463
FE9FF06F00078513
FFE7F79300052783
FD010113FE9FF06F
0291222302812423
0211262301312E23
01412C2303212023
0161282301512A23
0301041301712623
0005A2230005A783
0017F79300050993
0005278300F5A023
0407966300058493
0010079300B9A023
0005A78300F52423
00F5A0230017E793
02C12083FD040113
0241248302812403
01C1298302012903
01412A8301812A03
00C12B8301012B03
0000806703010113
00010A9300852783
0137879300279793
40F10133FF07F793
000A061300010A13
00251793A91FF0EF
FFC92B8300FA0933
00050B130049A783
00048513000B8593
00154593000780E7
000B851300048613
A3DFF0EF0FF5F593
001B0B130004A783
FFE7F79300992023
000B0B9300F4A023
0010081300090793
000A270301784A63
0017E79300072783
FFC7A6030CC0006F
00062703FFC78913
0A071E6300177713
FF878493FF87A583
000706930045A703
0005A68300E61663
04068063FFE6F693
000487930006A503
0205186300157513
FFEB8B930005A703
00E5A023FFE77713
0017671300062703
0006A70300E62023
00E6A02300176713
002B9793F81FF06F
FFC7A78300FA07B3
40E6073300462683
40D787B300173713
00F708630017B793
000A0513000B8593
FFFB8593A19FF0EF
A0DFF0EF000A0513
000727830004A703
00F720230017E793
0007278300092703
00F72023FFE7F793
0167D4630089A783
000A27830169A423
000A811300F9A023
FD010113E61FF06F
0291222302812423
0161282301412C23
0181242301712623
0321202302112623
01512A2301312E23
0301041301912223
00010B9300852783
0027979300050B13
FF07F79301378793
00010A1340F10133
00058493000A0613
00251C138E1FF0EF
FFCC2783018A0C33
0004A90310979263
FFE9791300050993
0044A7830C090463
001007930C078063
0137D46300000513
012C2023FF8C2503
0049278300198713
0007099300271A93
0E079E63015A0AB3
10050263FF8AAC83
0009061300452583
0015B593409585B3
0F949A63851FF0EF
0004A78300092703
0017F793FFE77713
00F4A02300E7E7B3
0017F79300092783
00F9202300F4E7B3
00F922230044A783
FFCC2783FFCAA703
FEEC2E230004A223
0004A683FEFAAE23
FFE6F79300092703
00F7673300177713
0009278300E4A023
FFE7F7930016F693
00F9202300D7E7B3
FFE7F9130004A783
0044A90300091463
0B374C6300100713
0A090463012B2023
0017E79300092783
000B811300F92023
02C12083FD040113
0241248302812403
01C1298302012903
01412A8301812A03
00C12B8301012B03
00412C8300812C03
0000806703010113
0017071300FAA023
EE9FF06F00078913
F11FF06F012B2023
00048613004CA583
412585B3000C8513
F44FF0EF0015B593
000926830004A703
FFE6F69300177793
00F4A02300D7E7B3
FFE7771300092783
00E7E7B30017F793
000B2423EF5FF06F
00299A93F65FF06F
FF8AA503015A0AB3
0017F79302091863
0607946300048613
0000061300452583
0015B593409585B3
000A2783EE0FF0EF
F29FF06F00FB2023
0009061300452583
0015B593409585B3
0004A783EC0FF0EF
000788630017F793
0017F79300092783
0009278300079A63
00F920230017E793
FF2AAE23FBDFF06F
0009859300000613
8A9FF0EF000A0513
00052503FA5FF06F
0005166300058793
0000806700000513
FFF007130085A683
80DFF06F00E69463
002697130005A603
0007250300E60733
FE0514E300452503
00D585330045A583
00050C6300054503
00D7A423FFF68693
00008067FFC72503
0087A68300E7A423
00D05863FFF68713
0006C68300D586B3
00E7A423FE0684E3
00271713F80748E3
0007250300E60733
FF01011300008067
0005851300050793
0006861300060593
000780E700112623
0EC030EF439020EF
0000806700000513
00812423FF010113
0450051300050413
0091222300112623
000400E700058493
0520051300048593
00040313000400E7
00C1208300812403
0041248300048593
0101011305200513
0005A78300030067
00F5A02300178793
07C7A303000067B7
FB01011300030067
03312E2304812423
03512A2303412C23
0411262303612823
0521202304912223
0381242303712623
03A1202303912223
00050A1301B12E23
0006099300058A93
0010041300068B13
0007041300E05463
02000C1300100793
03000C1300FB1463
001009133B9AD4B7
0000071300A00C93
00200D939FF48493
00148B9300A00D13
0934F26300071463
000A85930379D533
0305051300190913
00100713000A00E7
00100793FFFC8C93
03A4D4B30379F9B3
000A8593FCFC96E3
000A00E703098513
4124043300300793
04C1208306FB0A63
0441248304812403
03C1298304012903
03412A8303812A03
02C12B8303012B03
02412C8302812C03
01C12D8302012D03
0000806705010113
F96DEAE3F9944CE3
000C0513000A8593
000A00E700E12623
00C1270300190913
000A8593F79FF06F
000A00E702000513
FE8048E3FFF40413
000067B7F8DFF06F
0000806706A7AE23
04812423FB010113
0521202304912223
03412C2303312E23
0391222303512A23
01B12E2303A12023
0361282304112623
0381242303712623
0005849300050413
00068D1300060A93
FFF0091300000A13
00000C9300000993
000AC50380000DB7
04C1208304051063
0441248304812403
03C1298304012903
03412A8303812A03
02C12B8303012B03
02412C8302812C03
01C12D8302012D03
0000806705010113
02500693000C9E63
0004859336D50A63
001A8A93000400E7
06400693FA5FF06F
06A6E26310D50E63
02A6EA6303900693
0ED5746303100693
34D50A6302D00693
0CF5006303000793
02E5126302500713
0250051300048593
15C0006F000400E7
1AD50E6305800693
2EE50E6306300713
0250051300048593
00048593000400E7
FD5FF06F000AC503
16D50A6307000693
0690069302A6E063
06C006930AD50263
0680069308D50A63
FC5FF06FF6D506E3
10D5066307500693
0730071302A6EE63
000D2C03FAE518E3
000C0B93004D0B13
26051863000BC503
00F9986300300793
41790BB3418B8BB3
000B0D1327704663
078006930C80006F
07A0069312D50463
00095E63FA9FF06F
FD05091328098863
00200993F00992E3
FE0948E3EFDFF06F
02D9093300A00693
01250933FD090913
001A0A13FE1FF06F
040A1263EDDFF06F
004D0D13000D2603
0004859302065063
00C1202302D00513
00012603000400E7
40C00633FFF90913
0009869300090713
0004051300048593
03C0006FC95FF0EF
FAEA0EE300100713
FF87F713007D0793
0047268300072603
01B6073300870D13
00D7073300C73733
00048593FA0700E3
BF5FF0EF00040513
E59FF06F00000C93
000D2603000A1863
F9DFF06F004D0D13
FEEA08E300100713
FF87F713007D0793
0007260300870D13
FC0710E300472703
FFF7C793800007B7
FB1FF06FF6C7F8E3
0300051300048593
00048593000400E7
000400E707800513
0010099300800913
0B46C26300100693
00012423000D2783
00F12223004D0D13
00000B9301000C13
0100089300012023
0081258300412503
002B1613FFF88B13
C3CFE0EF01112623
0805186300F57513
0300069300012783
00C1288300079863
08F8966300100793
0185151300A68533
4185551300048593
001B8B93000400E7
00300693040B1863
D6D998E300000C93
41770BB300191713
00048593F17054E3
000400E702000513
FEDFF06FFFFB8B93
FF87F693007D0793
00868D130006A783
0046A78300F12223
F55FF06F00F12423
000B089301912023
00900793F59FF06F
F8A7E2E305700693
F7DFF06F03000693
00F12623FFFC0793
0010079301894C63
0004859300F99C63
000400E703000513
FC1FF06F00C12C03
FEF99AE300200793
0200051300048593
00048593FE5FF06F
000400E7001B8B93
00048593D81FF06F
000400E702000513
D85FF06FFFFB8B93
00048593000D2503
000400E7004D0B13
00000A13D75FF06F
00000993FFF00913
C89FF06F00100C93
C81FF06F00300993
C79FF06F00100993
00050613FE010113
0005869300002537
00C105939D450513
0001262300112E23
01C12083BA1FF0EF
0000806702010113
02B12223FC010113
00112E2302410593
02D1262302C12423
02F12A2302E12823
03112E2303012C23
FA5FF0EF00B12623
0401011301C12083
000065B700008067
FF01011300006537
D0050513CEC58593
0011262301E00613
000065B7FA9FF0EF
0060051391058593
00008067A99FE0EF
3007A7F300800793
0000806710500073
00A7953300100793
0000806730452573
3007B7F300800793
3440507330405073
FF01011300008067
0091222300812423
0011262300006437
0005049300A00793
00F51C630F040413
00D0059300042503
0047A78300452783
00042503000780E7
004527830FF4F593
000780E70047A783
0081240300C12083
0041248300048513
0000806701010113
0545051300002537
00006537A75FF06F
D0C50513FF010113
574000EF00112623
0EA7A823000067B7
00C12083FD9FF0EF
0101011300000513
800017B700008067
0207A5030247A703
FEE59AE30247A583
FE01011300008067
00112E2300812C23
0121282300912A23
0141242301312623
0080041301512223
0000693730043473
008474130F490513
02051E6358C020EF
000065B7000064B7
D3C5859300006537
D204861304E00693
E4DFF0EFC9850513
D545051300006537
04E00593E41FF0EF
E71FF0EFD2048513
000064B70F490513
0D84849359C020EF
0004A983F65FF0EF
000507130044AA83
00A7373341350533
0003D637415585B3
0000069309060613
8F4FE0EF40E585B3
090787930003D7B7
00050A1302A787B3
013789B30F490513
015787B300F9B7B3
00F4A2230134A023
02051E6350C020EF
000065B7000064B7
D6C5859300006537
D204861306100693
DA5FF0EFC9850513
D845051300006537
06100593D99FF0EF
DC9FF0EFD2048513
0181240330042473
0141248301C12083
00C1298301012903
000A051300412A83
0201011300812A03
FF0101136DD0206F
E99FF0EF00112623
090787930003D7B7
00F507B380001737
02D72623FFF00693
00B5053300A7B533
02A7262302F72423
DA5FF0EF00700513
0000051300C12083
0000806701010113
FE01011316059C63
00812C2300112E23
0121282300912A23
FFF0079301312623
0000453700F51663
000047B731A50513
31A78793FFF50413
000784131287DA63
3004B4F300800493
0F49051300006937
3D8020EF0084F493
000069B702051E63
00006537000065B7
04E00693D3C58593
C9850513D2098613
00006537C99FF0EF
C8DFF0EFD5450513
D209851304E00593
0F490513CBDFF0EF
DB9FF0EF3EC020EF
000067B70003D6B7
0D87879309068613
0047A5830007A703
08F6869302C407B3
3E70069340E68433
00F507B3008787B3
40A7053302C7D7B3
00F5053302C787B3
00C787B300A6C463
00E78733800016B7
02C6A623FFF00613
00B787B300F737B3
02F6A62302E6A423
348020EF0F490513
0000643702051E63
00006537000065B7
06100693D6C58593
C9850513D2040613
00006537BE1FF0EF
BD5FF0EFD8450513
D204051306100593
3004A4F3C05FF0EF
0181240301C12083
0101290301412483
0201011300C12983
EC045AE300008067
ECDFF06F00000413
FF01011300008067
0011262300812423
0121202300912223
3004347300800413
0F49051300006937
288020EF00847413
000064B702051E63
00006537000065B7
04E00693D3C58593
C9850513D2048613
00006537B49FF0EF
B3DFF0EFD5450513
D204851304E00593
0F490513B6DFF0EF
C69FF0EF29C020EF
0D87A483000067B7
0003D537409504B3
02A4D4B309050513
248020EF0F490513
0000693702051E63
00006537000065B7
06100693D6C58593
C9850513D2090613
00006537AE1FF0EF
AD5FF0EFD8450513
D209051306100593
30042473B05FF0EF
0081240300C12083
0001290300048513
0101011300412483
0005478300008067
00E794630005C703
40E7853300079663
0015051300008067
FE1FF06F00158593
000507930FF5F693
040718630037F713
008597130FF5F593
0105971300B765B3
00C7833300B765B3
0030081300078713
03186E6340E308B3
0027159300265713
FFC0059300B787B3
00C7073302B70733
02E7946300E78733
FE060EE300008067
FED78FA300178793
F9DFF06FFFF60613
FEB72E2300470713
00178793FB9FF06F
FD1FF06FFED78FA3
0000806700000513
00008067FDD00513
0087A78300052783
00B780230007A783
0025171300008067
00150513000067B7
00251513DAC78793
00E78733FF010113
0081242300A787B3
0007240300912223
001126230007A483
00C1208300946C63
0041248300812403
0000806701010113
0004051300042783
000780E70047A783
0004222300050463
FCDFF06F00C40413
000067B7FF010113
000064B700912223
0011262300812423
0121202309478413
0C44849309478793
0005091300941C63
0294146300078413
0440006F00000413
0007086300442703
0007270300042703
00C4041302A70863
00442783FD1FF06F
00C4041300079663
00042783FCDFF06F
0007A58300090513
FE0514E3E4DFF0EF
00C1208300040513
0041248300812403
0101011300012903
FF01011300008067
0091222300812423
0080041300112623
300437F300200493
00A4C46304D020EF
0010059300100513
90DFF0EF119020EF
00006537FE5FF06F
0D850613000067B7
40C7863354478793
0D85051300000593
FF010113DF9FF06F
0011262300200513
00006537E95FF0EF
85DFF0EFDC050513
E81FF0EF00300513
9B0FE0EF220020EF
4A078793000067B7
FFE7771300C7C703
00C1208300E78623
0000806701010113
08812C23F6010113
00006437000087B7
5507879309312623
00F9A22351040993
0700061301010793
0007851300000593
08912A2308112E23
D6DFF0EF09212823
00A9A42300100713
00E10EA300000513
00100513E05FF0EF
10100793DFDFF0EF
1CD010EF00F11E23
E0478793000067B7
00F1222300006937
00100793000026B7
4A090493000075B7
0000071300F12023
0000089300000793
73C6869300000813
7505859340000613
0299A0234A090513
00D4C7835C9010EF
FFB7F71351040413
01B7F79300E486A3
0184A78300079A63
4A09051300079663
000067B7134010EF
00F12223E0C78793
0010079300006537
000085B7000026B7
00F1202343050493
0000081302800893
0000071300000793
200006136E468693
43050513B5058593
00D4C783559010EF
0080051300942623
00F486A3FFB7F793
52878793000067B7
00F42E2300F42C23
0085751330053573
000067B7951FD0EF
FF0101135107A703
0011262300812423
0007841300912223
000064B702070E63
00006537000065B7
10000693E8458593
C9850513E6048613
00006537E98FF0EF
E8CFF0EFE9C50513
E604851310000593
51040793EBCFF0EF
00F7C7030087A783
02F71E6300100793
000065B700006437
EA05859300006537
E604061310100693
E4CFF0EFC9850513
E9C5051300006537
10100593E40FF0EF
E70FF0EFE6040513
51078793000067B7
00F747830087A703
00F707A3FFF78793
0081240300C12083
0101011300412483
0005242300008067
00A5202300052623
0000806700A52223
02812423FD010113
0005041301412C23
0291222302112623
01312E2303212023
00058A1301512A23
00C42703EF5FF0EF
51078793000067B7
0084260302070063
04D60E630087A683
609000EF060A1063
0280006FFF000513
00E686830087A683
001707130087A783
00E4262300D42823
5E1000EF00F42423
02C1208300000513
0241248302812403
01C1298302012903
01412A8301812A03
0000806703010113
FBDFF06F01042683
00E6890300E60783
000789130127D463
0000091300095463
3009B9F300800993
0F848513000064B7
439010EF0089F993
00006AB702051E63
00006537000065B7
04E00693D3C58593
C9850513D20A8613
00006537CF8FF0EF
CECFF0EFD5450513
D20A851304E00593
0F848513D1CFF0EF
0084250344D010EF
00F9566300E50783
558010EF00090593
00040613000A0693
0F84851300098593
00A126234BC010EF
509000EF00051863
F29FF06F00C12503
0104298300042783
00078C6300F40E63
0137D46300E78783
0009D46300078993
0080091300000993
0F84851330093973
381010EF00897913
00006A3702051E63
00006537000065B7
04E00693D3C58593
C9850513D20A0613
00006537C40FF0EF
C34FF0EFD5450513
D20A051304E00593
0F848513C64FF0EF
00842503395010EF
00F9866300E50783
4A0010EF00098593
349010EF0F848513
0000643702051E63
00006537000065B7
06100693D6C58593
C9850513D2040613
00006537BE0FF0EF
BD4FF0EFD8450513
D204051306100593
30092973C04FF0EF
FF500513425000EF
00C52783E45FF06F
00812C23FE010113
00912A2300112E23
0131262301212823
02079E6300050413
000065B7000064B7
E285859300006537
E14486130D400693
B74FF0EFC9850513
E9C5051300006537
0D400593B68FF0EF
B98FF0EFE1448513
00842703000067B7
02F70E635187A783
000065B7000064B7
E405859300006537
E14486130D500693
B2CFF0EFC9850513
E9C5051300006537
0D500593B20FF0EF
B50FF0EFE1448513
00C42783C3DFF0EF
02E7846300100713
00F42623FFF78793
01C1208301812403
0101290301412483
0201011300C12983
008004933450006F
000069373004B4F3
0084F4930F890513
02051E631E5010EF
000065B7000069B7
D3C5859300006537
D209861304E00693
AA4FF0EFC9850513
D545051300006537
04E00593A98FF0EF
AC8FF0EFD2098513
1F9010EF0F890513
0104258300842503
00F5846300E50783
00040513304010EF
00A424236C0000EF
06050A6300050993
01F7F79300D54783
0185278300079863
429000EF00079463
181010EF0F890513
0000693702051E63
00006537000065B7
06100693D6C58593
C9850513D2090613
00006537A18FF0EF
A0CFF0EFD8450513
D209051306100593
3004A4F3A3CFF0EF
0609A62300E98783
EF5FF06F00F42823
0F89051300042623
02051E63125010EF
000065B700006437
D6C5859300006537
D204061306100693
9BCFF0EFC9850513
D845051300006537
061005939B0FF0EF
9E0FF0EFD2040513
EA5FF06F3004A4F3
01F7F79300D54783
0185250300079863
0000806700153513
0000806700000513
00E5868300E50703
00D74C6300100793
00E6C86300000793
0105A50301052783
0007851300A7B7B3
FF01011300008067
DB0FF0EF00112623
1047A783000067B7
0000673700C12083
52A7202300A78533
0007851300000593
1940206F01010113
FF01011300052783
0011262300812423
0005041300912223
000064B702079863
00006537000065B7
C9850513F0458593
EF04861318300693
183005938E0FF0EF
910FF0EFEF048513
00C1208300042503
0041248300812403
0000806701010113
00812C23FE010113
0141242301212823
00912A2300112E23
0005091301312623
0080041300058A13
000064B730043473
008474130FC48513
02051E6379C010EF
000065B7000069B7
D3C5859300006537
D209861304E00693
85CFF0EFC9850513
D545051300006537
04E00593850FF0EF
880FF0EFD2098513
7B0010EF0FC48513
5207A023000067B7
00A0079300990913
000067B702F94933
000067B71127A223
EC9FF0EF1147A023
750010EF0FC48513
000064B702051E63
00006537000065B7
06100693D6C58593
C9850513D2048613
00006537FE9FE0EF
FDDFE0EFD8450513
D204851306100593
3004247380CFF0EF
0181240301C12083
0101290301412483
00812A0300C12983
0000806702010113
00812C23FE010113
00112E2301212823
0131262300912A23
0080041300050913
000064B730043473
008474130FC48513
02051E63694010EF
000065B7000069B7
D3C5859300006537
D209861304E00693
F55FE0EFC9850513
D545051300006537
04E00593F49FE0EF
F79FE0EFD2098513
6A8010EF0FC48513
E15FF0EF00890513
2F0000EF00090593
0FC4851300D94783
00F906A3FFD7F793
02051E63654010EF
000065B7000064B7
D6C5859300006537
D204861306100693
EEDFE0EFC9850513
D845051300006537
06100593EE1FE0EF
F11FE0EFD2048513
01C1208330042473
0009242301812403
0101290301412483
0201011300C12983
000067B700008067
FF0101135107A783
0011262300812423
0005841300912223
5D0010EF04079E63
000064B702051E63
00006537000065B7
07800693D6C58593
C9850513D2048613
00006537E69FE0EF
E5DFE0EFD8450513
D204851307800593
00040513E8DFE0EF
00C1208300812403
0101011300412483
578010EF8B0FD06F
000064B702051E63
00006537000065B7
06100693D6C58593
C9850513D2048613
00006537E11FE0EF
E05FE0EFD8450513
D204851306100593
00847413E35FE0EF
00C1208330042473
0041248300812403
0000806701010113
5107270300006737
844FD06F00071463
3007A7F300857793
0080051300008067
0085751330053573
FE010113FD9FF06F
00112E2300812C23
0121282300912A23
0080041301312623
000064B730043473
008474130FC48513
02051E6349C010EF
000065B700006937
D3C5859300006537
D209061304E00693
D5DFE0EFC9850513
D545051300006537
04E00593D51FE0EF
D81FE0EFD2090513
000069370FC48513
510927834AC010EF
02078E6351090913
000065B7000069B7
E845859300006537
E609861310000693
D0DFE0EFC9850513
E9C5051300006537
10000593D01FE0EF
D31FE0EFE6098513
00F7C70300892783
02F71E6300100793
000065B7000069B7
EA05859300006537
E609861310100693
CC5FE0EFC9850513
E9C5051300006537
10100593CB9FE0EF
CE9FE0EFE6098513
00F7478300892703
00F707A3FFF78793
3D8010EF0FC48513
000064B702051E63
00006537000065B7
06100693D6C58593
C9850513D2048613
00006537C71FE0EF
C65FE0EFD8450513
D204851306100593
30042473C95FE0EF
0181240301C12083
0101290301412483
0201011300C12983
000067B700008067
FF0101130907A783
0011262300812423
0005841300912223
000064B702F59863
00006537000065B7
C9850513F4858593
EF04861328C00693
28C00593BF9FE0EF
C29FE0EFEF048513
0004278300442703
0041248300C12083
00E7A22300F72023
0004222300042023
0101011300812403
0005278300008067
0000079300F51463
0000806700078513
01212823FE010113
00112E2301312623
00912A2300812C23
0080091300050993
000064B730093973
008979130FC48513
02051E63294010EF
000065B700006437
D3C5859300006537
D204061304E00693
B55FE0EFC9850513
D545051300006537
04E00593B49FE0EF
B79FE0EFD2040513
2A8010EF0FC48513
F71FF0EF00098513
0FC4851300050413
02051E63264010EF
000065B7000069B7
D6C5859300006537
D209861306100693
AFDFE0EFC9850513
D845051300006537
06100593AF1FE0EF
B21FE0EFD2098513
0C04066330092973
3009397300800913
008979130FC48513
02051E631E4010EF
000065B7000069B7
D3C5859300006537
D209861304E00693
AA5FE0EFC9850513
D545051300006537
04E00593A99FE0EF
AC9FE0EFD2098513
1F8010EF0FC48513
965FF0EF00840513
E41FF0EF00040593
0FC4851300D44783
00F406A3FFD7F793
02051E631A4010EF
000065B7000064B7
D6C5859300006537
D204861306100693
A3DFE0EFC9850513
D845051300006537
06100593A31FE0EF
A61FE0EFD2048513
0004242330092973
0B9010EF01840513
01C1208300040513
0141248301812403
00C1298301012903
0000806702010113
02812423FD010113
0321202302912223
01312E2302112623
000067B703010413
000504930907A783
02F5986300058913
000065B7000069B7
F485859300006537
2B000693C9850513
9A5FE0EFEF098613
EF0985132B000593
00C4A7039D5FE0EF
00F4A62300170793
04079A6300E92823
002797130084A783
FF07771301770713
40E1013301778793
00F10713FF07F793
00F1079340F10133
FF077713FF07F793
FFF00793FCF42C23
FCF42E23FCE42A23
00048513FD440593
02051863A54FE0EF
0004851300090593
FD040113D9DFD0EF
0281240302C12083
0201290302412483
0301011301C12983
00C4A78300008067
00E4A62300178713
FB5FF06F00F52823
0907A783000067B7
00812423FF010113
0011262300912223
0005041301212023
02F5986300058493
000065B700006937
F485859300006537
2CB00693C9850513
8ADFE0EFEF090613
EF0905132CB00593
000485938DDFE0EF
F11FD0EF00040513
0007946300042783
00C1208300042623
0041248300812403
0101011300012903
0000059300008067
FF010113CB1FD06F
0000643700812423
0005091301212023
0245051351040513
0011262300912223
51040413FD5FF0EF
0005146300050493
06091E6300C42483
02079E6300842783
000065B700006937
F1C5859300006537
EF09061307F00693
805FE0EFC9850513
E9C5051300006537
07F00593FF8FE0EF
829FE0EFEF090513
00D7C70300842783
0207166301F77713
07F0071300E7D683
02F4202302D77063
0081240300C12083
0001290300412483
0000806701010113
0097846300842783
02942023E5CFF0EF
FE010113FD9FF06F
0000693701212823
0087A78351090793
00812C2300112E23
00912A2300F7C783
5109091301312623
0000643702079E63
00006537000065B7
22100693EC858593
C9850513EF040613
00006537F50FE0EF
F44FE0EFE9C50513
EF04051322100593
00092783F74FE0EF
0000643702078E63
00006537000065B7
22200693E8458593
C9850513EF040613
00006537F10FE0EF
F04FE0EFE9C50513
EF04051322200593
00800413F34FE0EF
000064B730043473
008474130FC48513
02051E635FD000EF
000065B7000069B7
D3C5859300006537
D209861304E00693
EBCFE0EFC9850513
D545051300006537
04E00593EB0FE0EF
EE0FE0EFD2098513
611000EF0FC48513
0010051300892703
0017879300F74783
E21FF0EF00F707A3
5C1000EF0FC48513
000064B702051E63
00006537000065B7
06100693D6C58593
C9850513D2048613
00006537E58FE0EF
E4CFE0EFD8450513
D204851306100593
30042473E7CFE0EF
01C1208301812403
0101290301412483
0201011300C12983
FE010113865FF06F
0121282300812C23
00912A2300112E23
0005091301312623
3004347300800413
0FC48513000064B7
509000EF00847413
000069B702051E63
00006537000065B7
04E00693D3C58593
C9850513D2098613
00006537DC8FE0EF
DBCFE0EFD5450513
D209851304E00593
0FC48513DECFE0EF
0000653751D000EF
5345051300090593
00D94783BA9FF0EF
0407E79300000513
D21FF0EF00F906A3
4C1000EF0FC48513
000064B702051E63
00006537000065B7
06100693D6C58593
C9850513D2048613
00006537D58FE0EF
D4CFE0EFD8450513
D204851306100593
30042473D7CFE0EF
0181240301C12083
0101290301412483
0201011300C12983
FF05278300008067
00812C23FE010113
00112E2301312623
0121282300912A23
0005041301412423
0C078463FE850993
3004B4F300800493
0FC9051300006937
3F9000EF0084F493
00006A3702051E63
00006537000065B7
04E00693D3C58593
C9850513D20A0613
00006537CB8FE0EF
CACFE0EFD5450513
D20A051304E00593
0FC90513CDCFE0EF
FF04051340D000EF
00098593B78FF0EF
FF544783855FF0EF
FFD7F7930FC90513
3B9000EFFEF40AA3
0000693702051E63
00006537000065B7
06100693D6C58593
C9850513D2090613
00006537C50FE0EF
C44FE0EFD8450513
D209051306100593
3004A4F3C74FE0EF
FF544783FE042823
FEB7F79300098513
A84FF0EFFEF40AA3
0181240302050463
0141248301C12083
00812A0301012903
00C1298300098513
DD9FF06F02010113
0181240301C12083
0101290301412483
00812A0300C12983
0000806702010113
00812C23FE010113
00112E2301312623
0121282300912A23
0005099301412423
3004347300800413
0FC48513000064B7
2B9000EF00847413
0000693702051E63
00006537000065B7
04E00693D3C58593
C9850513D2090613
00006537B78FE0EF
B6CFE0EFD5450513
D209051304E00593
00006937B9CFE0EF
510909130FC48513
02490A132C5000EF
000A051300098593
00098593A51FF0EF
945FF0EF000A0513
0089250300D9C783
413505330407E793
00F986A300153513
0FC48513AB5FF0EF
02051E63255000EF
000065B7000064B7
D6C5859300006537
D204861306100693
AECFE0EFC9850513
D845051300006537
06100593AE0FE0EF
B10FE0EFD2048513
01C1208330042473
0141248301812403
00C1298301012903
0201011300812A03
000067B700008067
060786631047A783
51078793000067B7
07F006930087A703
04C6EA6300E75603
00E70603000066B7
04D642631006A683
0906A683000066B7
0187268302D70C63
0107A68302069863
FF01011302D54063
0011262300070513
00C12083E81FF0EF
8F8FF06F01010113
00D7A82340A686B3
FE01011300008067
0131262300812C23
00912A2300112E23
0005099301212823
3004347300800413
0FC48513000064B7
121000EF00847413
0000693702051E63
00006537000065B7
04E00693D3C58593
C9850513D2090613
000065379E0FE0EF
9D4FE0EFD5450513
D209051304E00593
0FC48513A04FE0EF
00D9C783135000EF
5109091300006937
00078E630407F793
0249051300098593
00D9C7838B1FF0EF
00F986A3FBF7F793
4135053300892503
921FF0EF00153513
0C1000EF0FC48513
000064B702051E63
00006537000065B7
06100693D6C58593
C9850513D2048613
00006537958FE0EF
94CFE0EFD8450513
D204851306100593
3004247397CFE0EF
0181240301C12083
0101290301412483
0201011300C12983
FE01011300008067
00912A2300812C23
0121282300050413
0131262300112E23
0006091300058493
00D44783EC5FF0EF
00F406A30027E793
000067B706048663
009424230907A783
000069B702F41863
00006537000065B7
C9850513F4858593
EF09861327600693
276005938B8FE0EF
8E8FE0EFEF098513
06F48C630004A783
00E4070306078A63
04D75C6300E78683
00F420230047A703
0087202300E42223
FFF007930087A223
0099091306F90463
02C9463300A00613
0181240301840513
0141248301C12083
00C1298301012903
A9458593000045B7
0016061302010113
0044A6834B90006F
0007A78300D78663
0044A783F8079CE3
00F4222300942023
0087A0230044A783
F99FF06F0084A223
0181240301C12083
0101290301412483
0201011300C12983
FF01011300008067
00812423000067B7
5187A50300050413
0005849300912223
0006861300060593
EB1FF0EF00112623
708000EF00040513
0000643702051E63
00006537000065B7
07800693D6C58593
C9850513D2040613
00006537FA1FD0EF
F95FD0EFD8450513
D204051307800593
00812403FC5FD0EF
0004851300C12083
0101011300412483
FE0101139E8FC06F
0121282300812C23
00112E2301312623
0141242300912A23
0005091301512223
0080041300058993
000064B730043473
008474130FC48513
02051E6364C000EF
000065B700006A37
D3C5859300006537
D20A061304E00693
F0DFD0EFC9850513
D545051300006537
04E00593F01FD0EF
F31FD0EFD20A0513
660000EF0FC48513
D4DFE0EF00090513
00050A9301899993
0A0508634189D993
534A0A1300006A37
000A051300090593
000A0513DD0FF0EF
0009059301390723
00100513CC0FF0EF
0FC48513E44FF0EF
02051E635E4000EF
000065B7000064B7
D6C5859300006537
D204861306100693
E7DFD0EFC9850513
D845051300006537
06100593E71FD0EF
EA1FD0EFD2048513
040A806330042473
5187A783000067B7
0207986300F7C783
01C1208301812403
0101290301412483
00812A0300C12983
0201011300412A83
0139072386CFF06F
01C12083F7DFF06F
0141248301812403
00C1298301012903
00412A8300812A03
0000806702010113
00003737000067B7
E387071351078793
0000051300000593
0207A6230207A223
02E7A4230207A823
00E50503D19FE06F
FE01011300008067
0000643700812C23
00112E2351042783
0121282300912A23
5104041301312623
000064B702078E63
00006537000065B7
37E00693E8458593
C9850513EF048613
00006537D81FD0EF
D75FD0EFE9C50513
EF04851337E00593
000067B7DA5FD0EF
0907A78300842703
008007930CF70663
000064B73007B7F3
0087F9930FC48513
02051E6345C000EF
000065B700006937
D3C5859300006537
D209061304E00693
D1DFD0EFC9850513
D545051300006537
04E00593D11FD0EF
D41FD0EFD2090513
470000EF0FC48513
0244091300842583
BFCFF0EF00090513
0009051300842583
00100513AF0FF0EF
0FC48513C74FF0EF
02051E63414000EF
000065B700006437
D6C5859300006537
D204061306100693
CADFD0EFC9850513
D845051300006537
06100593CA1FD0EF
CD1FD0EFD2040513
008005133009A7F3
0181240330053573
0141248301C12083
00C1298301012903
0201011300857513
FD010113EE1FB06F
000064B702912223
028124235104A783
0321202302112623
01412C2301312E23
5104849300050413
0000693702078E63
00006537000065B7
39800693E8458593
C9850513EF090613
00006537C19FD0EF
C0DFD0EFE9C50513
EF09051339800593
02041663C3DFD0EF
00040513E35FF0EF
0281240302C12083
0201290302412483
01812A0301C12983
0000806703010113
001409930AC010EF
0001262300A98433
3009397300800913
0089791300C10513
02051E632CC000EF
000065B700006A37
D3C5859300006537
D20A061304E00693
B8DFD0EFC9850513
D545051300006537
04E00593B81FD0EF
BB1FD0EFD20A0513
2E0000EF00C10513
931FF0EF0084A503
000045B70084A503
0185051300098613
7C4000EFA9458593
00C105130084A703
0107E79300D74783
278000EF00F706A3
000069B702051E63
00006537000065B7
07800693D6C58593
C9850513D2098613
00006537B11FD0EF
B05FD0EFD8450513
D209851307800593
00090513B35FD0EF
0084A783D69FB0EF
0107F79300D7C783
000064B702078E63
00006537000065B7
3B500693F5C58593
C9850513EF048613
00006537AC1FD0EF
AB5FD0EFE9C50513
EF0485133B500593
781000EFAE5FD0EF
EA0454E340A40433
EA1FF06F00000413
00812423FF010113
0091222300112623
00050413FFF00793
000064B702F51E63
00006537000065B7
3C400693F3C58593
C9850513EF048613
00006537A59FD0EF
A4DFD0EFE9C50513
EF0485133C400593
00940413A7DFD0EF
02A4453300A00513
3E800793DCDFF0EF
0640061302F515B3
02F5053300000693
00C12083D19FB0EF
0041248300812403
0000806701010113
5187A503000067B7
00D5478300008067
0007986301F7F793
0015351301852503
0000051300008067
000067B700008067
00A035335107A503
000067B700008067
00C7C5035187A783
0000806700157513
02012303FE010113
00112E2300812C23
0005041300612023
000067B7E8CFC0EF
01C120835187A783
06F424230687A783
0201011301812403
0605278300008067
00812423FF010113
0005041300112623
000780E700078463
F61FF0EF00040513
0004051302050463
00D44783F14FF0EF
0087E79300C12083
0081240300F406A3
0000806701010113
0027F79300D44783
0004051300078663
01842783971FE0EF
01840513FC0786E3
FC1FF06F7AC000EF
00C506A300D50623
000507A300B50723
00052E2300052C23
0005250300008067
000067B700050E63
003575135247C783
00A0353340F50533
0010051300008067
000067B700008067
0147C70351078793
00E7E7B30087A783
00F7186300052703
0010051300052023
0000051300008067
000067B700008067
0147C70351078793
00E7E7B30087A783
0000806700F52023
00812C23FE010113
00112E2301212823
0131262300912A23
0080041300050913
000064B730043473
0084741310848513
02051E63F5DFF0EF
000065B7000069B7
D3C5859300006537
D209861304E00693
81DFD0EFC9850513
D545051300006537
04E00593811FD0EF
841FD0EFD2098513
F71FF0EF10848513
0047F71300D94783
1084851306071463
02051E63F2DFF0EF
000065B7000064B7
D6C5859300006537
D204861306100693
FC4FD0EFC9850513
D845051300006537
06100593FB8FD0EF
FE8FD0EFD2048513
01C1208330042473
0141248301812403
00C1298301012903
0000806702010113
00F906A3FFB7F793
D89FF0EF00090513
0009051300050663
00040593954FF0EF
01C1208301812403
00C1298301012903
0141248310848513
8A1FE06F02010113
03512223FC010113
000066B700068A93
02812C235106A683
0331262302912A23
02112E2303412423
0005049303212823
00060A1300058993
04068E6304412403
000065B700006937
1B30069300006537
E8458593F9490613
01112E23C9850513
00F12A2301012C23
EDCFD0EF00E12823
FA85051300006537
1B300593ED0FD0EF
F00FD0EFF9490513
0181280301C12883
0101270301412783
0001222304012683
00D12023000A0613
000A869300098593
CE5FF0EF00048513
00F40863FFF00793
0004851302041A63
03C12083E11FF0EF
0004851303812403
0341248303012903
02812A0302C12983
0401011302412A83
0094041300008067
02C4463300A00613
A9458593000045B7
0016061301848513
FB9FF06F2B0000EF
000067B7FD010113
0000693703212023
0291222302812423
01312E2302112623
0C47841301412C23
0C4909130C478493
0004841303246E63
FFF0049384DFE0EF
00004A3700A00993
0281240307246463
0241248302C12083
01C1298302012903
0301011301812A03
02C42783E2DFE06F
0204278300F12223
0144278300F12023
0184280301C42883
00C4268301042703
0044258300842603
BE5FF0EF00042503
0487AE2300042783
F85FF06F03040413
0096086302442603
0006186300042503
03040413D01FF0EF
00960613F81FF06F
A94A059303364633
0016061301850513
FE1FF06F1C8000EF
00812C23FE010113
00112E2300912A23
0005049301212823
0080041300012623
00C1051330043473
C39FF0EF00847413
0000693702051E63
00006537000065B7
04E00693D3C58593
C9850513D2090613
00006537CF8FD0EF
CECFD0EFD5450513
D209051304E00593
00C10513D1CFD0EF
00C4C783C4DFF0EF
02078E630017F793
000065B700006937
FE85859300006537
FD09061302900693
CACFD0EFC9850513
01C5051300006537
02900593CA0FD0EF
CD0FD0EFFD090513
B19FF0EF00048513
00C1051300040593
01C12083DD4FE0EF
0141248301812403
0201011301012903
000067B700008067
0007946310C7A783
000005138C5FD06F
0005278300008067
0000673702050263
00E50C6308472703
0087A70300078A63
00D7073300852683
0045270300E7A423
00E7A22300F72023
0005222300052023
000067B700008067
FF0101131147C783
0081242300112623
FFF0051300912223
8000053700079663
000067B7FFF54513
0007A40308078793
0204026302F40463
F69FF0EF00842483
0000051340A484B3
008424030004C863
40A40533F55FF0EF
5207A783000067B7
00A7D46300078663
00C1208300078513
0041248300812403
0000806701010113
FD01011300052783
0291222302812423
0211262301312E23
01412C2303212023
0161282301512A23
0181242301712623
0005899300050413
02078E6300060493
000065B700006937
04C5859300006537
0389061305400693
B2CFD0EFC9850513
E9C5051300006537
05400593B20FD0EF
B50FD0EF03890513
0090446301342623
0080099300100493
00006A373009B9F3
0089F993110A0513
02051E63A0DFF0EF
000065B700006937
D3C5859300006537
D209061304E00693
ACCFD0EFC9850513
D545051300006537
04E00593AC0FD0EF
AF0FD0EFD2090513
A21FF0EF110A0513
00950533E45FF0EF
0804A903000064B7
0804849300A42423
00006AB700990C63
00006BB700006B37
0209106300006C37
009420230044A783
0044A78300F42223
0084A2230087A023
0089278305C0006F
06CB05930207D663
038A861305D00693
A44FD0EFC98B8513
A3CFD0EFE9CC0513
038A851305D00593
00892703A6CFD0EF
0AE7D86300842783
00F9242340F707B3
0124202300492783
0087A02300F42223
0004A78300892223
00F4186300978A63
00000593DEDFF0EF
110A0513CE0FD0EF
02051E6392DFF0EF
000065B700006437
D6C5859300006537
D204061306100693
9C4FD0EFC9850513
D845051300006537
061005939B8FD0EF
9E8FD0EFD2040513
02C120833009A9F3
0241248302812403
01C1298302012903
01412A8301812A03
00C12B8301012B03
0301011300812C03
40E787B300008067
0044A78300F42423
00092903EF2788E3
FE010113EE5FF06F
0131262300812C23
00912A2300112E23
0005099301212823
3004347300800413
11048513000064B7
849FF0EF00847413
0000693702051E63
00006537000065B7
04E00693D3C58593
C9850513D2090613
00006537908FD0EF
8FCFD0EFD5450513
D209051304E00593
1104851392CFD0EF
0009A78385DFF0EF
00078863FEA00913
C89FF0EF00098513
1104851300000913
02051E6380DFF0EF
000065B7000064B7
D6C5859300006537
D204861306100693
8A4FD0EFC9850513
D845051300006537
06100593898FD0EF
8C8FD0EFD2048513
01C1208330042473
0009051301812403
0101290301412483
0201011300C12983
FF01011300008067
0011262300812423
0121202300912223
3004347300800413
11048513000064B7
F58FF0EF00847413
0000693702051E63
00006537000065B7
04E00693D3C58593
C9850513D2090613
00006537818FD0EF
80CFD0EFD5450513
D209051304E00593
1104851383CFD0EF
BE9FF0EFF6CFF0EF
1104851300050913
02051E63F2CFF0EF
000065B7000064B7
D6C5859300006537
D204861306100693
FC5FC0EFC9850513
D845051300006537
06100593FB9FC0EF
FE9FC0EFD2048513
00C1208330042473
0009051300812403
0001290300412483
0000806701010113
00812C23FE010113
0141242301212823
00912A2300112E23
0005091301312623
0080041300058A13
000064B730043473
0084741311048513
02051E63E6CFF0EF
000065B7000069B7
D3C5859300006537
D209861304E00693
F2DFC0EFC9850513
D545051300006537
04E00593F21FC0EF
F51FC0EFD2098513
E80FF0EF11048513
00A95C63AFDFF0EF
00A7D86300100793
00090513000A0593
110485139E0FD0EF
02051E63E2CFF0EF
000065B7000064B7
D6C5859300006537
D204861306100693
EC5FC0EFC9850513
D845051300006537
06100593EB9FC0EF
EE9FC0EFD2048513
01C1208330042473
0141248301812403
00C1298301012903
0201011300812A03
FD01011300008067
01412C2302812423
0291222302112623
01312E2303212023
0161282301512A23
0181242301712623
01A1202301912223
0080041300050A13
30043473B9DFE0EF
1109051300006937
D50FF0EF00847413
000064B702051E63
00006537000065B7
04E00693D3C58593
C9850513D2048613
00006537E11FC0EF
E05FC0EFD5450513
D204851304E00593
000069B7E35FC0EF
D60FF0EF11090513
1149A623000064B7
10C9899300006A37
0E048493080A0A13
00006BB700006AB7
00006C3700006B37
000A2D0300006CB7
0004A6830009A783
014D0C630044A503
008D2703000D0A63
40F707330AE7DC63
00D786B300ED2423
00A7073341F7D713
00E787B300F6B7B3
00F4A22300D4A023
969FF0EF0009A023
85CFD0EF00000593
CA8FF0EF11090513
000064B702051E63
00006537000065B7
06100693D6C58593
C9850513D2048613
00006537D41FC0EF
D35FC0EFD8450513
D204851306100593
30042473D65FC0EF
0281240302C12083
0201290302412483
01812A0301C12983
01012B0301412A83
00812C0300C12B83
00012D0300412C83
0000806703010113
41F7559300D706B3
00E6B63300A585B3
40E787B300B60633
000D2423000D0513
00C4A22300D4A023
871FF0EF00F9A023
BF8FF0EF11090513
D6CB859302051663
D20A861306100693
C9DFC0EFC98B0513
C95FC0EFD84C0513
D20A851306100593
30042473CC5FC0EF
000D051300CD2783
000780E700800413
1109051330043473
B80FF0EF00847413
D3CC859302051863
D20A861304E00693
C4DFC0EFC98B0513
D545051300006537
04E00593C41FC0EF
C71FC0EFD20A8513
BA0FF0EF11090513
FE010113E6DFF06F
00112E2300912A23
0121282300812C23
0080049301312623
000069373004B4F3
0084F49311090513
02051E63B14FF0EF
000065B700006437
D3C5859300006537
D204061304E00693
BD5FC0EFC9850513
D545051300006537
04E00593BC9FC0EF
BF9FC0EFD2040513
B28FF0EF11090513
000067B781CFD0EF
0007A9830E078793
013509B30047A403
0085043300A9B533
AD0FF0EF11090513
0000693702051E63
00006537000065B7
06100693D6C58593
C9850513D2090613
00006537B69FC0EF
B5DFC0EFD8450513
D209051306100593
3004A4F3B8DFC0EF
01C1208300040593
0009851301812403
0101290301412483
0201011300C12983
FF01011300008067
EF9FF0EF00112623
0101011300C12083
FF01011300008067
FE1FF0EF00112623
02F535B33E800793
0000069306400613
DEDFA0EF02F50533
0101011300C12083
FF01011300008067
0091222300812423
000064B700006437
0C44041300112623
00946E630C448493
0081240300C12083
0000051300412483
0000806701010113
0004051301440793
00F42C2300F42A23
01C40413929FB0EF
00008067FCDFF06F
00000C1C00000000
00000C1C00000000
00000C1C00000000
00000C1C00000000
00000C1C00000000
00000C1C00000000
00000C1C00000000
0000210C00000000
000020C40000590C
00005D1400000000
0000000000002254
000025B800005D0C
0000590C00006088
00000000000054D4
0303030302020100
0404040404040404
0505050505050505
0505050505050505
0606060606060606
0606060606060606
0606060606060606
0606060606060606
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0000612C00006118
0000615400006140
0000617C00006168
007365786574756D
0063696D616E7964
35315B1B4A325B1B
206F6D654448313B
7470697263736544
2D2D2D2D0A6E6F69
2D2D2D2D2D2D2D2D
206E410A2D2D2D2D
6E656D656C706D69
6F206E6F69746174
756C6F7320612066
206F74206E6F6974
696E694420656874
6F6C69685020676E
0A73726568706F73
206D656C626F7270
7373616C63206128
69746C756D206369
206461657268742D
6E6F7268636E7973
206E6F6974617A69
296D656C626F7270
7020736968540A2E
616C756369747261
6D656C706D692072
6E6F697461746E65
74736E6F6D656420
6874207365746172
2065676173752065
69746C756D20666F
656572700A656C70
20656C626974706D
706F6F6320646E61
2065766974617265
2073646165726874
656666696420666F
69727020676E6972
2C7365697469726F
6C6C65770A736120
2520732520736120
687420646E612073
656C732064616572
000A2E676E697065
5320202020202020
20474E4956524154
0000202020202020
49444C4F48202020
4620454E4F20474E
00002020204B524F
474E495441452020
64257325205B2020
0000205D20736D20
50504F5244202020
4620454E4F204445
00002020204B524F
4E494B4E49485420
64257325205B2047
0000205D20736D20
0000005000000043
4864253B64255B1B
6C69685000000000
20726568706F736F
253A73255B206425
000000205D642573
00000BAC00000AF4
00000AE800000BAC
00000B9400000AF4
0000596000000BA0
0000599C00005980
000059BC000059B0
6E6B6E75000059D4
65637845006E776F
6163206E6F697470
2820732520657375
000000000A296425
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
7463757274736E49
72646461206E6F69
6173696D20737365
000064656E67696C
7463757274736E49
65636341206E6F69
746C756166207373
656C6C4900000000
74736E69206C6167
006E6F6974637572
696F706B61657242
64616F4C0000746E
7373657264646120
67696C6173696D20
64616F4C0064656E
2073736563636120
000000746C756166
72654B202A2A2A2A
6F6C6C41206C656E
46206E6F69746163
20216572756C6961
0000000A2A2A2A2A
654B202A2A2A2A2A
504F4F206C656E72
2A2A2A2A2A202153
2A2A2A2A0000000A
6C656E72654B202A
202163696E615020
00000A2A2A2A2A2A
6B6E55202A2A2A2A
746146206E776F6E
726F727245206C61
2A2A2A2021642520
7272754300000A2A
6572687420746E65
203D204449206461
746C7561460A7025
74736E6920676E69
206E6F6974637572
2073736572646461
200A78257830203D
257830203A617220
30203A7067202078
3A70742020782578
7420207825783020
0A78257830203A30
7830203A31742020
203A327420207825
3374202078257830
202078257830203A
78257830203A3474
30203A357420200A
3A36742020782578
6120207825783020
2078257830203A30
257830203A316120
203A326120200A78
3361202078257830
202078257830203A
78257830203A3461
7830203A35612020
3A366120200A7825
6120207825783020
0A78257830203A37
0052534900000000
6169746E65737365
646165726874206C
6174614600000000
20746C756166206C
5320217325206E69
2E676E696E6E6970
61746146000A2E2E
20746C756166206C
6165726874206E69
6241202170252064
0A2E676E6974726F
7275705300000000
746E692073756F69
6420747075727265
2164657463657465
6425203A51524920
72612F2E0000000A
76637369722F6863
2F65726F632F3233
632E646165726874
2828282800000000
797469726F697270
3034203D3D202929
73695F7A20262620
68745F656C64695F
6874282864616572
6E75665F64616572
207C7C2029292963
202D203034282828
2828203D3E202931
262029292939322D
6F69727028282026
3E20292979746972
2939322D2828203D
7028282026262029
29797469726F6972
303428203D3C2029
0029292931202D20
4F49545245535341
5B204C494146204E
73252040205D7325
000000000A64253A
64696C61766E6909
7469726F69727020
203B296425282079
206465776F6C6C61
25203A65676E6172
0A6425206F742064
696C2F2E00000000
7373612F736F2F62
000000632E747265
3A64253A73252040
747261750000000A
5F73797300000030
0000006B636F6C63
2E2E2F2E2E2F2E2E
6564756C636E692F
636F6C6E6970732F
70735F7A00682E6B
5F6B636F6C5F6E69
296C2864696C6176
6365520900000000
7320657669737275
0A6B636F6C6E6970
70735F7A00000000
636F6C6E755F6E69
2864696C61765F6B
746F4E090000296C
6E69707320796D20
00000A216B636F6C
000025C8000025C0
0000000000000000
0000609400000000
000060C4000060B8
000060C4000060C4
6F42202A2A2A2A2A
655A20676E69746F
20534F2072796870
762D72796870657A
312D302E34312E31
333331672D303331
3231623037383736
0A2A2A2A2A2A2032
6E69616D00000000
656C646900000000
656B2F2E00000000
74756D2F6C656E72
00000000632E7865
6C3E2D786574756D
6E756F635F6B636F
00005530203E2074
6F3E2D786574756D
203D3D2072656E77
2E6C656E72656B5F
00746E6572727563
2E2E2F2E2E2F2E2E
2F6C656E72656B2F
2F6564756C636E69
682E64656863736B
6B5F282100000000
656E2E6C656E7265
203D212064657473
00000A0900295530
2E6C656E72656B5F
2D746E6572727563
63732E657361623E
6B636F6C5F646568
0031203D21206465
2E6C656E72656B5F
2D746E6572727563
63732E657361623E
6B636F6C5F646568
0030203D21206465
6C656E72656B2F2E
632E64656863732F
6572687400000000
657361623E2D6461
5F6465646E65702E
72656B5F00006E6F
727275632E6C656E
28203D2120746E65
292A2064696F7628
2120736D00002930
000029312D28203D
656C64695F736921
2964616572687428
695F7A2100000000
6461657268745F73
735F65746174735F
6E72656B5F287465
65727275632E6C65
55312828202C746E
293428203C3C204C
656B2F2E00292929
7268742F6C656E72
000000632E646165
7364616572685409
746F6E2079616D20
6165726320656220
49206E6920646574
000000000A735253
6C656E72656B2F2E
5F6461657268742F
00632E74726F6261
2D64616572687428
73752E657361623E
6F6974706F5F7265
312828202620736E
3028203C3C204C55
203D3D2029292929
7373650900005530
74206C6169746E65
6261206461657268
00000A646574726F
6C656E72656B2F2E
74756F656D69742F
737973210000632E
695F65646F6E645F
64656B6E696C5F73
6F6E3E2D6F742628
643E2D7400296564
3D3E20736B636974
0000198000003020
0000608000006080
FFFFFFF580001008
0000559400006430
0000000000000000
00005D9800005588
0000557000000000
0000000000000000
000000000000557C
000060C400000000
00000000000060C4
0000002800000000
