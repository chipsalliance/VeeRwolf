@00000000
37 05 00 10 13 05 05 00 B7 05 00 00 93 85 05 03 
83 82 05 00 23 00 55 00 93 85 15 00 83 82 05 00 
E3 9A 02 FE B7 05 00 20 93 85 05 00 23 A0 05 00 
@00000030
53 77 65 52 56 2B 46 75 73 65 53 6F 43 20 72 6F 
63 6B 73 0A 00 
