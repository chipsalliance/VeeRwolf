0102829300000297
13D0006F30529073
00112023FB010113
0041242300312223
0061282300512623
01C12C2300712A23
03E1202301D12E23
02A1242303F12223
02C1282302B12623
02E12C2302D12A23
0501202302F12E23
341022F305112223
300022F304512423
1F0000EF04512623
02051E6300000313
800003B7342022F3
0072F2B3FFF38393
00628A6300B00313
0000009700010513
7E40006F13408093
0042829304812283
0900006F04512423
0000339700010293
0043A103B3838393
00512023FF010113
001E0E130003AE03
0003086301C3A023
03C0809300000097
3420257302D0006F
FFF28293800002B7
158000EF00557533
4302829300002297
00A282B300351513
0042A3030002A503
00003317000300E7
00032383AD830313
00732023FFF38393
0002811300012283
02032E0300832383
00003297087E0863
0082A303AB028293
0293282302832623
03332C2303232A23
0553202303432E23
0573242305632223
0593282305832623
05B32C2305A32A23
0000339702232423
0003AE0391838393
0202A30307C32623
028321030062A423
0303248302C32403
0383298303432903
04032A8303C32A03
04832B8304432B03
05032C8304C32C03
05832D8305432D03
3412907304812283
3002907304C12283
0041218300012083
00C1228300812203
0141238301012303
01C12E8301812E03
02412F8302012F03
02C1258302812503
0341268303012603
03C1278303812703
0441288304012803
3020007305010113
0000329700000073
0082A3039C028293
0085751306C32383
00038513300522F3
0010031300008067
3442B37300A312B3
342022F300008067
0062F2B380000337
0002846300000513
0000806700150513
0200079302060063
00F04C6340C787B3
00000713FE060513
0007059300A5D533
00C5D73300008067
00F595B300C55533
FE9FF06F00B56533
0006081300058793
0005031300068893
0000273728069663
0EC5F66359870713
0CD67863000106B7
00C6B6B30FF00693
00D658B300369693
0007470301170733
0200071300D706B3
00070C6340D70733
00D556B300E797B3
00F6E5B300E61833
0108551300E51333
0108161302A5F733
0103569301065613
0107171302A5D5B3
02B607B300D766B3
00F6FE6300058713
FFF58713010686B3
00F6F6630106E863
010686B3FFE58713
02A6F7B340F686B3
0103531301031313
0107979302A6D6B3
02D605B30067E333
00B37C6300068513
FFF6851300680333
00B3746301036663
01071713FFE68513
0000059300A76733
010008B70E40006F
F3166CE301000693
F31FF06F01800693
0010069300061663
000106B702C6D833
0FF006930CD87263
008008930106F463
00D70733011856B3
0200071300074683
40D70733011686B3
410787B30A071863
0108561300100593
0108D89301081893
02C7F73301035693
0107171302C7D7B3
02F8853300D766B3
00A6FE6300078713
FFF78713010686B3
00A6F6630106E863
010686B3FFE78713
02C6F7B340A686B3
0103531301031313
0107979302C6D6B3
02D888B30067E333
01137C6300068513
FFF6851300680333
0113746301036663
01071713FFE68513
0007051300A76733
010006B700008067
F4D862E301000893
F3DFF06F01800893
00D7D5B300E81833
00D556B300E51333
00E797B301085513
00F6E8B302A5F733
0107D79301081793
02A5D5B30108D613
00C7673301071713
0005861302B786B3
0107073300D77E63
01076863FFF58613
FFE5861300D77663
40D706B301070733
0108989302A6F733
02A6D6B30108D893
02D785B301071713
00068713011767B3
010787B300B7FE63
0107E863FFF68713
FFE6871300B7F663
40B787B3010787B3
00E5E5B301061593
18D5E663EB5FF06F
04E6F46300010737
00D837330FF00813
0000283700371713
00E6D5B359880813
0005C803010585B3
00E8083302000593
02059663410585B3
EEF6ECE300100713
0015471300C53533
010005B7EEDFF06F
FCB6E0E301000713
FB9FF06F01800713
00B696B301065733
0106DE9300D766B3
03D778B30107D733
0105583300B797B3
0106979300F86333
010358130107D793
03D7573300B61633
0108E83301089893
00070E1302E78F33
00D8083301E87E63
00D86863FFF70E13
FFE70E1301E87663
41E8083300D80833
03D8583303D878B3
03078EB301089893
0107D79301031793
0008071300F8E7B3
00D787B301D7FE63
00D7E863FFF80713
FFE8071301D7F663
010E1E1300D787B3
00010EB741D787B3
FFFE881300EE6733
0107589301077333
0106561301067833
0308883303030E33
02C30333010E5693
006686B301030333
0106F46302C888B3
0106D61301D888B3
0317E663011608B3
000107B7CF179AE3
00F6F6B3FFF78793
00FE7E3301069693
01C686B300B51533
DAD57CE300000593
CC9FF06FFFF70713
0000071300000593
000025B7DA5FF06F
6985859300002537
2DD0006F6A850513
00112623FF010113
0060079300812423
75C010EF02F50463
754010EF02050463
000035B704051663
0000353796C58593
2A5000EF98050513
FFDFF06F2E1000EF
FC051CE3740010EF
BEC4041300003437
0000353700842583
27D000EF9A050513
161010EF00842503
000035B7FD1FF06F
FB9FF06F96858593
04812423FB010113
0411262304912223
0005049300600793
0EA7E06300058413
0025179300002737
00E787B36BC70713
000780670007A783
7EC5051300002537
688010EF221000EF
0104288304442783
02F1282300C42803
0044270304042783
02F1262300042683
0484260303C42783
02F1242300050593
0000353703842783
02F1222387050513
02F1202303442783
00F12E2303042783
00F12C2302C42783
00F12A2302842783
00F1282302442783
00F1262302042783
00F1242301C42783
00F1222301842783
00F1202301442783
18D000EF00842783
0004851300040593
00003537EA9FF0EF
F55FF06F81450513
8305051300003537
00003537F49FF06F
84C5051300048593
F39FF06F159000EF
00812423FF010113
0005041300112623
0016161334202673
0050079300165613
0000273702C7E863
6D87071300261793
0007A58300F707B3
6F85051300002537
00040593111000EF
EA5FF0EF00000513
6F058593000025B7
FF010113FE1FF06F
342025F300112623
0015959300003537
9C8505130015D593
000025B70D9000EF
0040051371458593
000037B7E69FF0EF
0007A703AF078793
0007A30300070C63
000037B70007A023
00030067AF47A503
FF01011300008067
5D9000EF00112623
63D000EF0F1000EF
8D81011300003117
80028293000012B7
FD9FF0EF00510133
FD01011321C0006F
0006899301312E23
0281242303012683
0005841303212023
0008859300060913
0291222300400613
0005049302112623
00F1242300E12623
6FC010EF01012223
FB09059300812783
0404AE2300B405B3
FF05F5930604A023
000027B702F5A823
0041280300C12703
04F5A62388078793
02C12083000017B7
9607879302812403
02E5A6230335A423
04F5A4230305AA23
0201290302B4A423
01C1298302412483
0000806703010113
02F5873300C00793
00E787B300C52783
00B7546300B50703
020007130007A783
01F6751302E64733
00E787B300271713
0000806700F6A023
00C10693FE010113
FBDFF0EF00112E23
0010079300C12703
0007278300A79533
00A7E7B301C12083
0201011300F72023
0045278300008067
FF01011300855803
02F8083300812423
0005250300050413
FFF0071300A44883
0091222300112623
0000059300E405A3
0105053300C00313
02000E9301F00E13
000004930315C263
06F4C46300845783
0081240300C12083
0101011300412483
02F8573300008067
026586B300C42603
0046861300D606B3
00C6A42300C6A223
00B405A300EE4E63
003787930027D793
00158593FFC7F793
01F70713FA9FF06F
00A6A02303D74733
00E5053300271713
00442783FD9FF06F
0000059300048613
0004278302F48733
0014849300040513
00C4270300E787B3
00D7A02300470693
00D7A22300872683
00F6A02300872683
ED5FF0EF00F72423
FF010113F51FF06F
0005851300050793
0006861300060593
000780E700112623
520010EF2A4010EF
0000806700000513
00812423FF010113
0450051300050413
0091222300112623
000400E700058493
0520051300048593
00040313000400E7
00C1208300812403
0041248300048593
0101011305200513
0005A78300030067
00F5A02300178793
A807A303000037B7
FB01011300030067
03312E2304812423
03512A2303412C23
0411262303612823
0521202304912223
0381242303712623
03A1202303912223
00050A1301B12E23
0006099300058A93
0010041300068B13
0007041300E05463
02000C1300100793
03000C1300FB1463
001009133B9AD4B7
0000071300A00C93
00200D939FF48493
00148B9300A00D13
0934F26300071463
000A85930379D533
0305051300190913
00100713000A00E7
00100793FFFC8C93
03A4D4B30379F9B3
000A8593FCFC96E3
000A00E703098513
4124043300300793
04C1208306FB0A63
0441248304812403
03C1298304012903
03412A8303812A03
02C12B8303012B03
02412C8302812C03
01C12D8302012D03
0000806705010113
F96DEAE3F9944CE3
000C0513000A8593
000A00E700E12623
00C1270300190913
000A8593F79FF06F
000A00E702000513
FE8048E3FFF40413
000037B7F8DFF06F
00008067A8A7A023
04812423FB010113
0521202304912223
03412C2303312E23
0391222303512A23
01B12E2303A12023
0361282304112623
0381242303712623
0005849300050413
00068D1300060A93
FFF0091300000A13
00000C9300000993
000AC50380000DB7
04C1208304051063
0441248304812403
03C1298304012903
03412A8303812A03
02C12B8303012B03
02412C8302812C03
01C12D8302012D03
0000806705010113
02500693000C9E63
0004859336D50A63
001A8A93000400E7
06400693FA5FF06F
06A6E26310D50E63
02A6EA6303900693
0ED5746303100693
34D50A6302D00693
0CF5006303000793
02E5126302500713
0250051300048593
15C0006F000400E7
1AD50E6305800693
2EE50E6306300713
0250051300048593
00048593000400E7
FD5FF06F000AC503
16D50A6307000693
0690069302A6E063
06C006930AD50263
0680069308D50A63
FC5FF06FF6D506E3
10D5066307500693
0730071302A6EE63
000D2C03FAE518E3
000C0B93004D0B13
26051863000BC503
00F9986300300793
41790BB3418B8BB3
000B0D1327704663
078006930C80006F
07A0069312D50463
00095E63FA9FF06F
FD05091328098863
00200993F00992E3
FE0948E3EFDFF06F
02D9093300A00693
01250933FD090913
001A0A13FE1FF06F
040A1263EDDFF06F
004D0D13000D2603
0004859302065063
00C1202302D00513
00012603000400E7
40C00633FFF90913
0009869300090713
0004051300048593
03C0006FC95FF0EF
FAEA0EE300100713
FF87F713007D0793
0047268300072603
01B6073300870D13
00D7073300C73733
00048593FA0700E3
BF5FF0EF00040513
E59FF06F00000C93
000D2603000A1863
F9DFF06F004D0D13
FEEA08E300100713
FF87F713007D0793
0007260300870D13
FC0710E300472703
FFF7C793800007B7
FB1FF06FF6C7F8E3
0300051300048593
00048593000400E7
000400E707800513
0010099300800913
0B46C26300100693
00012423000D2783
00F12223004D0D13
00000B9301000C13
0100089300012023
0081258300412503
002B1613FFF88B13
A1CFF0EF01112623
0805186300F57513
0300069300012783
00C1288300079863
08F8966300100793
0185151300A68533
4185551300048593
001B8B93000400E7
00300693040B1863
D6D998E300000C93
41770BB300191713
00048593F17054E3
000400E702000513
FEDFF06FFFFB8B93
FF87F693007D0793
00868D130006A783
0046A78300F12223
F55FF06F00F12423
000B089301912023
00900793F59FF06F
F8A7E2E305700693
F7DFF06F03000693
00F12623FFFC0793
0010079301894C63
0004859300F99C63
000400E703000513
FC1FF06F00C12C03
FEF99AE300200793
0200051300048593
00048593FE5FF06F
000400E7001B8B93
00048593D81FF06F
000400E702000513
D85FF06FFFFB8B93
00048593000D2503
000400E7004D0B13
00000A13D75FF06F
00000993FFF00913
C89FF06F00100C93
C81FF06F00300993
C79FF06F00100993
00050613FE010113
0005869300001537
00C10593BF450513
0001262300112E23
01C12083BA1FF0EF
0000806702010113
02B12223FC010113
00112E2302410593
02D1262302C12423
02F12A2302E12823
03112E2303012C23
FA5FF0EF00B12623
0401011301C12083
0000806700008067
3007A7F300800793
0000806710500073
00A7953300100793
0000806730452573
3007B7F300800793
3440507330405073
FF01011300008067
0091222300812423
0011262300003437
0005049300A00793
00F51C63AF840413
00D0059300042503
0047A78300452783
00042503000780E7
004527830FF4F593
000780E70047A783
0081240300C12083
0041248300048513
0000806701010113
00812423FF010113
2444051300001437
320000EF00112623
0081240324440513
0101011300C12083
00003537A85FF06F
9F050513FF010113
394000EF00112623
AEA7AC23000037B7
00C12083FB9FF0EF
0101011300000513
800017B700008067
0207A5030247A703
FEE59AE30247A583
FE01011300008067
00112E2300812C23
0121282300912A23
0080041301312623
000034B730043473
FC1FF0EFAE048493
0044A9830004A903
4125053300050713
413585B300A73733
090606130003D637
40E585B300000693
0003D7B7F41FE0EF
02A787B309078793
0127893300847413
013787B300F937B3
00F4A2230124A023
0181240330042473
0141248301C12083
00C1298301012903
7C50006F02010113
00112623FF010113
0003D7B7F45FF0EF
8000173709078793
FFF0069300F507B3
00A7B53302D72623
02F7242300B50533
0070051302A72623
00C12083E31FF0EF
0101011300000513
0C059C6300008067
00812423FF010113
0091222300112623
00050413FFF00793
000047B700F51663
0080049331A78413
ED1FF0EF3004B4F3
FFF4079300004737
0084F49331A70713
0007079308F75463
090705930003D737
000037B702B786B3
0007A603AE078793
08F707930047A803
00A787B340C787B3
3E70071340A60533
02B7D7B300D787B3
00F5053302B787B3
00B787B300A74463
00C7863380001737
02D72623FFF00693
010787B300F637B3
02F7262302C72423
00C120833004A4F3
0041248300812403
0000806701010113
00000793F807D0E3
00008067F79FF06F
00812423FF010113
0080041300112623
E11FF0EF30043473
AE07A783000037B7
40F5053300847413
090787930003D7B7
3004247302F55533
0081240300C12083
0000806701010113
0005C70300054783
0007966300E79463
0000806740E78533
0015859300150513
0FF5F693FE1FF06F
0037F71300050793
0FF5F59304071863
00B765B300859713
00B765B301059713
0007871300C78333
40E308B300300813
0026571303186E63
00B787B300271593
02B70733FFC00593
00E7873300C70733
0000806702E79463
00178793FE060EE3
FFF60613FED78FA3
00470713F9DFF06F
FB9FF06FFEB72E23
FED78FA300178793
FFF00513FD1FF06F
000037B700008067
00008067A8A7A223
0000806700000513
00008067FDD00513
0087A78300052783
00B780230007A783
0025171300008067
00150513000037B7
00251513A1878793
00E78733FF010113
0081242300A787B3
0007240300912223
001126230007A483
00C1208300946C63
0041248300812403
0000806701010113
0004051300042783
000780E70047A783
0004222300050463
FCDFF06F00C40413
000037B7FF010113
000034B700912223
0011262300812423
01212023A9C78413
ACC48493A9C78793
0005091300941C63
0294146300078413
0440006F00000413
0007086300442703
0007270300042703
00C4041302A70863
00442783FD1FF06F
00C4041300079663
00042783FCDFF06F
0007A58300090513
FE0514E3E39FF0EF
00C1208300040513
0041248300812403
0101011300012903
0000353700008067
AE050613000037B7
40C78633C1878793
AE05051300000593
FF010113E1DFF06F
0011262300200513
00003537ECDFF0EF
A85FF0EFA2C50513
EB9FF0EF00300513
F89FE0EF061000EF
B7C78793000037B7
FFE7771300C7C703
00C1208300E78623
0000806701010113
08812C23F6010113
00003437000047B7
A207879309312623
00F9A223BEC40993
0700061301010793
0007851300000593
08912A2308112E23
D91FF0EF09212823
00A9A42300100713
00E10EA300000513
00100513E3DFF0EF
10100793E35FF0EF
638000EF00F11E23
A7078793000037B7
00F1222300003937
00100793000016B7
B7C90493000035B7
0000071300F12023
0000089300000793
7346869300000813
C205859340000613
0299A023B7C90513
00D4C7836D8000EF
FFB7F713BEC40413
01B7F79300E486A3
0184A78300079A63
B7C9051300079663
000037B72DC000EF
00F12223A7878793
0010079300003537
000035B7000026B7
00F12023B0C50493
0000081300F00893
0000071300000793
2000061349468693
B0C5051302058593
00D4C783668000EF
0080051300942623
00F486A3FFB7F793
C0478793000037B7
00F42E2300F42C23
0085751330053573
00452703959FE0EF
00F7202300052783
0005202300E7A223
0000806700052223
01F7F79300D54783
0185250300079863
0000806700153513
0000806700000513
00112623FF010113
000037B7BC9FF0EF
00C12083B007A783
00A7853300003737
00000593BEA72E23
0101011300078513
FF0101131E10006F
0011262300812423
3004347300800413
BE07AE23000037B7
00A0079300950513
000037B702F54533
B0A7A02300847413
AEB7AE23000037B7
30042473F91FF0EF
0081240300C12083
0000806701010113
00812423FF010113
0011262300912223
0080041300050493
F21FF0EF30043473
0084741300D4C783
00F486A3FFD7F793
00C1208330042473
0004A42300812403
0101011300412483
000037B700008067
00079663BEC7A783
835FE06F00058513
3005A5F30085F593
0000373700008067
00071463BEC72703
00857793819FE06F
000080673007A7F3
3005357300800513
FD9FF06F00857513
3007B7F300800793
BF47268300003737
FFF7071300F6C703
0087F79300E687A3
000080673007A7F3
00F5146300052783
0007851300000793
FE01011300008067
0000343700812C23
0005049300912A23
02450513BEC40513
FCDFF0EF00112E23
00051463BEC40413
0084278300C42503
00D7C70302049A63
0207146301F77713
07F0071300E7D683
02F4202300D77E63
0181240301C12083
0201011301412483
00F5086300008067
E35FF0EF00A12623
02A4202300C12503
FF010113FD9FF06F
0011262300812423
3004347300800413
BF47A703000037B7
0084741300100513
0017879300F74783
F51FF0EF00F707A3
0081240330042473
0101011300C12083
FF010113EF1FF06F
0011262300812423
3004347300800413
BEC7079300003737
000036B70247A783
00847413C1068693
06D78063BEC70713
0287258304078E63
00E7880300E50603
0047A70305065063
00E5222300F52023
00A7A22300A72023
0407E79300D54783
0000051300F506A3
30042473ECDFF0EF
0081240300C12083
0000806701010113
0007A78300B78663
02872783FA079AE3
00F5222300D52023
00A7A02302872783
FB5FF06F02A72423
FF010113FF052783
0121202300812423
0091222300112623
FE85091300050413
0080049302078663
000905133004B4F3
FF544783CC5FF0EF
FFD7F7930084F493
3004A4F3FEF40AA3
FF544783FE042823
FEB7F79300090513
CB5FF0EFFEF40AA3
0081240302050063
0041248300C12083
0001290300090513
ED9FF06F01010113
0081240300C12083
0001290300412483
0000806701010113
00812423FF010113
0011262300912223
0080049300050413
C41FF0EF3004B4F3
BEC7079300003737
000036B70247A783
0084F493C1068693
06D78663BEC70713
0287258306078463
00E7850300E40603
0047A68304A65663
00D4222300F42023
0087A2230086A023
0087250300D44783
408505330407E793
0015351300F406A3
3004A4F3D75FF0EF
0081240300C12083
0101011300412483
00B7866300008067
FA0794E30007A783
00D4202302872783
0287278300F42223
028724230087A023
000037B7FA9FF06F
06078663B007A783
BEC78793000037B7
07F006930087A703
04C6EA6300E75603
00E70603000036B7
04D64263AFC6A683
A986A683000036B7
0187268302D70C63
0107A68302069863
FF01011302D54063
0011262300070513
00C12083EE1FF0EF
B6DFF06F01010113
00D7A82340A686B3
FF01011300008067
0091222300812423
0005049300112623
3004347300800413
0084741300D54783
00078A630407F793
00D4C783AF5FF0EF
00F486A3FBF7F793
BF47A503000037B7
0015351340950533
30042473C6DFF0EF
0081240300C12083
0101011300412483
000037B700008067
02478713BEC78793
02E7A42302E7A223
0000051300000593
000037B7B0DFF06F
00008067BF47A503
01F7F79300D54783
0185250300079863
0000806700153513
0000806700000513
BEC7A503000037B7
0000806700A03533
BF47A783000037B7
0015751300C7C503
FF01011300008067
0011262300812423
0080041300912223
00D5478330043473
0047F71300847413
3004247300071E63
0081240300C12083
0101011300412483
FFB7F79300008067
0005049300F506A3
00050663F71FF0EF
C51FF0EF00048513
0081240300040593
0041248300C12083
C185051300003537
AE1FF06F01010113
02012303FE010113
00112E2300812C23
0005041300612023
000037B7A45FE0EF
01C12083BF47A783
06F424230687A783
0201011301812403
0605278300008067
00812423FF010113
0005041300112623
000780E700078463
EE5FF0EF00040513
0004051302050463
00D44783E45FF0EF
0087E79300C12083
0081240300F406A3
0000806701010113
0027F79300D44783
0004051300078663
018427839F9FF0EF
01840513FC0786E3
FC1FF06F2FC000EF
000037B7FD010113
0000393703212023
0291222302812423
01312E2302112623
ACC7841301412C23
ACC90913ACC78493
0004841303246E63
FFF00493A41FF0EF
00002A3700A00993
0281240307246463
0241248302C12083
01C1298302012903
0301011301812A03
02C42783ACDFF06F
0204278300F12223
0144278300F12023
0184280301C42883
00C4268301042703
0044258300842603
EB5FF0EF00042503
0487AE2300042783
F85FF06F03040413
0096086302442603
0006186300042503
03040413E15FF0EF
00960613F81FF06F
BE0A059303364633
0016061301850513
FE1FF06F134000EF
00C506A300D50623
000507A300B50723
00052E2300052C23
FD01011300008067
0080059302112623
0085F5933005B5F3
E71FF0EF00B12623
01C1051300C12583
02C12083905FF0EF
0000806703010113
B047A783000037B7
BE4FF06F00079463
0000806700000513
0205026300052783
A8C7270300003737
00078A6300E50C63
008526830087A703
00E7A42300D70733
00F7202300452703
0005202300E7A223
0000806700052223
B087C783000037B7
00112623FF010113
0091222300812423
00079663FFF00513
FFF5451380000537
A8878793000037B7
02F404630007A403
0084248302040263
40A484B3F69FF0EF
0004C86300000513
F55FF0EF00842403
000037B740A40533
00078663BFC7A783
0007851300A7D463
0081240300C12083
0101011300412483
FE01011300008067
00912A2300812C23
0005041300112E23
00B5262300C12623
3004B4F300800493
00C12603F01FF0EF
00C044630084F493
000037B700100613
00A60633A887A703
A887879300C42423
0047A58300F70663
0047A70302071063
00E4222300F42023
008720230047A703
02C0006F0087A223
0084268300872603
40D606B304C6D863
0047268300D72423
00D4222300E42023
008722230086A023
00F70A630007A703
ED5FF0EF00E41863
988FF0EF00000593
01C120833004A4F3
0141248301812403
0000806702010113
00D4242340C686B3
00072703F8B702E3
FF010113F79FF06F
0011262300812423
3004347300800413
0084741300052783
E3DFF0EF02078063
3004247300000513
0081240300C12083
0000806701010113
FE9FF06FFEA00513
00112623FF010113
0080079300812423
E45FF0EF3007B473
3007A7F300847793
0081240300C12083
0000806701010113
00812C23FE010113
00112E2300912A23
00B1262300050493
3004347300800413
00847413E09FF0EF
00A4DA6300C12583
00A7D66300100793
8A8FF0EF00048513
01C1208330042473
0141248301812403
0000806702010113
00812C23FE010113
00112E2300912A23
0131262301212823
0151222301412423
0080041300050493
3004347399DFF0EF
00003A37000039B7
B099A22300003937
B049899300847413
AE890913A88A0A13
000A248300800A93
000926830009A783
01448C6300492503
0084A70300048A63
40F7073306E7D063
00D786B300E4A423
00A7073341F7D713
00E787B300F6B7B3
00F9222300D92023
D35FF0EF0009A023
FE9FE0EF00000593
01C1208330042473
0141248301812403
00C1298301012903
00412A8300812A03
0000806702010113
41F7559300D706B3
00E6B63300A585B3
40E787B300B60633
000485130004A423
00C9222300D92023
C95FF0EF00F9A023
00C4A78330042473
000780E700048513
00847413300AB473
FF010113F3DFF06F
0091222300812423
0080041300112623
300437F300200493
00A4C463E41FF0EF
0010059300100513
D4DFE0EFE61FF0EF
FF010113FE5FF06F
0091222300812423
000034B700003437
ACC4041300112623
00946E63ACC48493
0081240300C12083
0000051300412483
0000806701010113
0004051301440793
00F42C2300F42A23
01C40413D64FE0EF
00008067FCDFF06F
000008DC00000000
000008DC00000000
000008DC00000000
000008DC00000000
000008DC00000000
000008DC00000000
000008DC00000000
0000131C00000000
000012D400002710
000029F800000000
00000000000013B8
000015E8000029F0
0000271000002A90
00000000000024CC
0303030302020100
0404040404040404
0505050505050505
0505050505050505
0606060606060606
0606060606060606
0606060606060606
0606060606060606
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
666C6F7672657773
0000737978656E5F
6F57206F6C6C6548
0A73252021646C72
000007B400000000
0000086C0000086C
000007B4000007A8
0000086000000854
0000278400002764
000027B4000027A0
000027D8000027C0
006E776F6E6B6E75
6F69747065637845
206573756163206E
0A29642528207325
DEADBAAD00000000
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
74736E49DEADBAAD
206E6F6974637572
2073736572646461
6E67696C6173696D
74736E4900006465
206E6F6974637572
6620737365636341
00000000746C7561
206C6167656C6C49
7463757274736E69
61657242006E6F69
0000746E696F706B
6464612064616F4C
73696D2073736572
0064656E67696C61
6363612064616F4C
6C75616620737365
2A2A2A2A00000074
206C656E72654B20
697461636F6C6C41
756C696146206E6F
2A2A2A2A20216572
2A2A2A2A0000000A
6C656E72654B202A
2A202153504F4F20
0000000A2A2A2A2A
654B202A2A2A2A2A
6E6150206C656E72
2A2A2A2A20216369
2A2A2A2A00000A2A
6E776F6E6B6E5520
45206C6174614620
21642520726F7272
00000A2A2A2A2A20
20746E6572727543
4920646165726874
460A7025203D2044
20676E69746C7561
7463757274736E69
72646461206E6F69
7830203D20737365
3A617220200A7825
6720207825783020
2078257830203A70
257830203A707420
30203A3074202078
317420200A782578
202078257830203A
78257830203A3274
7830203A33742020
203A347420207825
7420200A78257830
2078257830203A35
257830203A367420
30203A3061202078
3A31612020782578
20200A7825783020
78257830203A3261
7830203A33612020
203A346120207825
3561202078257830
200A78257830203A
257830203A366120
30203A3761202078
000000000A782578
6573736500525349
6874206C6169746E
0000000064616572
6166206C61746146
25206E6920746C75
6E6E697053202173
000A2E2E2E676E69
6166206C61746146
74206E6920746C75
7025206461657268
6974726F62412021
000000000A2E676E
73756F6972757053
75727265746E6920
6365746564207470
5152492021646574
0000000A6425203A
0000003074726175
636F6C635F737973
000015F00000006B
00000000000015F8
0000000000000000
00002AC000002A9C
00002ACC00002ACC
2A2A2A2A00002ACC
6E69746F6F42202A
72796870655A2067
6870657A20534F20
34312E31762D7279
2D303331312D302E
3738373633333167
2A2A203232316230
000000000A2A2A2A
000000006E69616D
00000000656C6469
000015D400000BA0
00002A8800002A88
FFFFFFF580001008
0000258C00002B0C
0000000000000000
00002A0400002580
0000256800000000
0000000000000000
0000000000002574
00002ACC00000000
0000000000002ACC
0000000F00000000
