0102829300000297
47D0006F30529073
00112023FB010113
0041242300312223
0061282300512623
01C12C2300712A23
03E1202301D12E23
02A1242303F12223
02C1282302B12623
02E12C2302D12A23
0501202302F12E23
341022F305112223
300022F304512423
1F0000EF04512623
02051E6300000313
800003B7342022F3
0072F2B3FFF38393
00628A6300B00313
0000009700010513
3250006F13408093
0042829304812283
0900006F04512423
0000639700010293
0043A10306838393
00512023FF010113
001E0E130003AE03
0003086301C3A023
03C0809300000097
3420257336D0006F
FFF28293800002B7
158000EF00557533
F882829300005297
00A282B300351513
0042A3030002A503
00006317000300E7
0003238300830313
00732023FFF38393
0002811300012283
02032E0300832383
00006297087E0863
0082A303FE028293
0293282302832623
03332C2303232A23
0553202303432E23
0573242305632223
0593282305832623
05B32C2305A32A23
0000639702232423
0003AE03B2438393
0202A30307C32623
028321030062A423
0303248302C32403
0383298303432903
04032A8303C32A03
04832B8304432B03
05032C8304C32C03
05832D8305432D03
3412907304812283
3002907304C12283
0041218300012083
00C1228300812203
0141238301012303
01C12E8301812E03
02412F8302012F03
02C1258302812503
0341268303012603
03C1278303812703
0441288304012803
3020007305010113
0000629700000073
0082A303EF028293
0085751306C32383
00038513300522F3
0010031300008067
3442B37300A312B3
342022F300008067
0062F2B380000337
0002846300000513
0000806700150513
0200079302060063
00F04C6340C787B3
00000713FE060513
0007059300A5D533
00C5D73300008067
00F595B300C55533
FE9FF06F00B56533
0006081300058793
0005031300068893
0000573728069663
0EC5F6630F070713
0CD67863000106B7
00C6B6B30FF00693
00D658B300369693
0007470301170733
0200071300D706B3
00070C6340D70733
00D556B300E797B3
00F6E5B300E61833
0108551300E51333
0108161302A5F733
0103569301065613
0107171302A5D5B3
02B607B300D766B3
00F6FE6300058713
FFF58713010686B3
00F6F6630106E863
010686B3FFE58713
02A6F7B340F686B3
0103531301031313
0107979302A6D6B3
02D605B30067E333
00B37C6300068513
FFF6851300680333
00B3746301036663
01071713FFE68513
0000059300A76733
010008B70E40006F
F3166CE301000693
F31FF06F01800693
0010069300061663
000106B702C6D833
0FF006930CD87263
008008930106F463
00D70733011856B3
0200071300074683
40D70733011686B3
410787B30A071863
0108561300100593
0108D89301081893
02C7F73301035693
0107171302C7D7B3
02F8853300D766B3
00A6FE6300078713
FFF78713010686B3
00A6F6630106E863
010686B3FFE78713
02C6F7B340A686B3
0103531301031313
0107979302C6D6B3
02D888B30067E333
01137C6300068513
FFF6851300680333
0113746301036663
01071713FFE68513
0007051300A76733
010006B700008067
F4D862E301000893
F3DFF06F01800893
00D7D5B300E81833
00D556B300E51333
00E797B301085513
00F6E8B302A5F733
0107D79301081793
02A5D5B30108D613
00C7673301071713
0005861302B786B3
0107073300D77E63
01076863FFF58613
FFE5861300D77663
40D706B301070733
0108989302A6F733
02A6D6B30108D893
02D785B301071713
00068713011767B3
010787B300B7FE63
0107E863FFF68713
FFE6871300B7F663
40B787B3010787B3
00E5E5B301061593
18D5E663EB5FF06F
04E6F46300010737
00D837330FF00813
0000583700371713
00E6D5B30F080813
0005C803010585B3
00E8083302000593
02059663410585B3
EEF6ECE300100713
0015471300C53533
010005B7EEDFF06F
FCB6E0E301000713
FB9FF06F01800713
00B696B301065733
0106DE9300D766B3
03D778B30107D733
0105583300B797B3
0106979300F86333
010358130107D793
03D7573300B61633
0108E83301089893
00070E1302E78F33
00D8083301E87E63
00D86863FFF70E13
FFE70E1301E87663
41E8083300D80833
03D8583303D878B3
03078EB301089893
0107D79301031793
0008071300F8E7B3
00D787B301D7FE63
00D7E863FFF80713
FFE8071301D7F663
010E1E1300D787B3
00010EB741D787B3
FFFE881300EE6733
0107589301077333
0106561301067833
0308883303030E33
02C30333010E5693
006686B301030333
0106F46302C888B3
0106D61301D888B3
0317E663011608B3
000107B7CF179AE3
00F6F6B3FFF78793
00FE7E3301069693
01C686B300B51533
DAD57CE300000593
CC9FF06FFFF70713
0000071300000593
FE010113DA5FF06F
00812C2300112E23
0006041300912A23
0121282300058493
305030EF00050913
00A1262375C030EF
0010061300005537
3E05051300190593
00C12703091010EF
0000563706074263
3DC60613000056B7
0000553740468693
3EC5051300090593
06040063069010EF
0487D6633E700793
45C58593000055B7
0004851300040613
01812403049010EF
0141248301C12083
0000553701012903
0201011355C50513
000056370290106F
3D860613000056B7
FA1FF06F45C68693
40458593000055B7
000055B7FB9FF06F
0004851345C58593
FB1FF06F7F8010EF
02912A23FC010113
02112E2303412423
0321282302812C23
0351222303312623
01712E2303612023
01912A2301812C23
01B1262301A12823
0005049300500793
0EF50E6300150A13
1F078793000057B7
00E7873300251713
002A171300072903
0007A98300E787B3
00005D3700005DB7
01900A9306400B13
00005C3700005CB7
0000061300005BB7
00048513360D8593
FFF00593E95FF0EF
5E5010EF00090513
378D059300000613
E79FF0EF00048513
00098513FFF00593
774040EF5C9010EF
390C859303655433
0344043300048513
0014041301F47413
0004061303540433
00040513E45FF0EF
00098513724030EF
3A8C05937CD010EF
0004851300000613
00090513E25FF0EF
724040EF7B5010EF
3C0B859303655433
0344043300048513
0014041301F47413
0004061303540433
00040513DF5FF0EF
F49FF06F6D4030EF
D249099300006937
D249091306498993
00005637F19FF06F
00005537000055B7
20860613FC010113
2185051321058593
02812C2302112E23
0321282302912A23
0341242303312623
0361202303512223
65C010EF01712E23
0000059300001537
214020EF38850513
D245041300006537
4B9010EFD2450513
4B1010EF01440513
4A9010EF02840513
4A1010EF03C40513
499010EF05040513
0000693706440513
489010EF00006437
15090913D9C40413
00300A9300000493
00400B13FFF00B93
0060099300000A37
00048713409A88B3
0000081300090593
7C0A069300000793
0004051330000613
0161202301712223
000405132D1030EF
19D030EF00148493
3009091307040413
03C12083FD3490E3
0341248303812403
02C1298303012903
02412A8302812A03
01C12B8302012B03
0000806704010113
00112623FF010113
0060079300812423
7E8030EF02F50463
7E0030EF02050463
000055B704051663
000055376B858593
544010EF6CC50513
FFDFF06F5B0010EF
FC051CE37CC030EF
11C4041300006437
0000553700842583
51C010EF6EC50513
425030EF00842503
000055B7FD1FF06F
FB9FF06F6B458593
04812423FB010113
0411262304912223
0005049300600793
0EA7E06300058413
0025179300005737
00E787B340870713
000780670007A783
5385051300005537
714030EF4C0010EF
0104288304442783
02F1282300C42803
0044270304042783
02F1262300042683
0484260303C42783
02F1242300050593
0000553703842783
02F122235BC50513
02F1202303442783
00F12E2303042783
00F12C2302C42783
00F12A2302842783
00F1282302442783
00F1262302042783
00F1242301C42783
00F1222301842783
00F1202301442783
42C010EF00842783
0004851300040593
00005537EA9FF0EF
F55FF06F56050513
57C5051300005537
00005537F49FF06F
5985051300048593
F39FF06F3F8010EF
00812423FF010113
0005041300112623
0016161334202673
0050079300165613
0000573702C7E863
4247071300261793
0007A58300F707B3
4445051300005537
000405933B0010EF
EA5FF0EF00000513
43C58593000055B7
FF010113FE1FF06F
342025F300112623
0015959300005537
714505130015D593
000055B7378010EF
0040051346058593
000067B7E69FF0EF
0007A703CF878793
0007A30300070C63
000067B70007A023
00030067CFC7A503
FF01011300008067
720010EF00112623
784010EF3D0010EF
CC81011300007117
80028293000012B7
FD9FF0EF00510133
FD0101134BD0006F
0291222302812423
01312E2303212023
01512A2301412C23
0171262301612823
0211262300078B13
0280079301812423
0005841300050493
00068A1300060993
00080A9300070B93
08F89A6300088913
36C78793000027B7
0301268308F69A63
0004851300090593
5F4030EF00400613
00B405B3FB098593
0404AE23000027B7
FF05F5930604A023
04F5A62388078793
02C12083000017B7
CA07879302812403
0375A6230345A423
0355AA230365A823
02B4A42304F5A423
0241248302012903
01812A0301C12983
01012B0301412A83
00812C0300C12B83
0000806703010113
0440079301D88693
00005C37F6D7FAE3
00006537000055B7
0180069373CC0613
8045051377858593
00006537200010EF
FE30069300090593
8245051302700613
018005931E8010EF
218010EF73CC0513
00C00793F2DFF06F
00C5278302F58733
00B5070300E787B3
0007A78300B75463
02E6473302000713
0027171301F67513
00F6A02300E787B3
FE01011300008067
00112E2300C10693
00C12703FBDFF0EF
00A7953300100793
01C1208300072783
00F7202300A7E7B3
0000806702010113
0085580300452783
00812423FF010113
0005041302F80833
00A4488300052503
00112623FFF00713
00E405A300912223
00C0031300000593
01F00E1301050533
0315C26302000E93
0084578300000493
00C1208306F4C463
0041248300812403
0000806701010113
00C4260302F85733
00D606B3026586B3
00C6A22300468613
00EE4E6300C6A423
0027D79300B405A3
FFC7F79300378793
FA9FF06F00158593
03D7473301F70713
0027171300A6A023
FD9FF06F00E50533
0004861300442783
02F4873300000593
0004051300042783
00E787B300148493
0047069300C42703
0087268300D7A023
0087268300D7A223
00F7242300F6A023
F51FF06FED5FF0EF
00C5222300058663
0005278300008067
00F666330017F793
0000806700C52023
FE01011300052783
00912A2300812C23
0131262301212823
0005099300112E23
00F6202300058913
0010049300060413
0325926300042583
0181240301C12083
0101290300048513
00C1298301412483
0000806702010113
000905130049A783
00042783000780E7
0047A78300051E63
FC0782E300440413
00F4202300148493
0007A783FB1FF06F
FE5FF06FFFE7F793
FD01011300259793
01612823FF878793
0321202300F50B33
00478793000B2903
00F504B302912223
0049278302812423
01412C230004A403
40F40A3301712623
01312E2302112623
001A3B9301512A23
00442A8308F41C63
08F40C6301403A33
0020079300442983
FFCB250300B7DE63
0045258300040613
0015B593412585B3
000A8613ED1FF0EF
00040513000B8593
00090613EC1FF0EF
00040513000A0593
00098613EB1FF0EF
00090513000B8593
02C12083EA1FF0EF
02812403008B2023
01C129830124A023
0201290302412483
01412A8301812A03
00C12B8301012B03
0000806703010113
FFEAFA9300042A83
00042983F69FF06F
F69FF06FFFE9F993
0005A7030085A783
0027969300178793
00D7073300F5A423
0045A70300A72023
00F707B300100693
0005250300078023
0005A7030085A783
00051A63FFE57513
00F707B300279793
000080670007A503
0027961300178793
00C7073300F5A423
0045A70300A72023
00D7802300F707B3
FD010113FBDFF06F
40000BB701712623
0161282301312E23
01A1202301812423
0281242302112623
0321202302912223
01512A2301412C23
00050D1301912223
00060B1300058993
FFFB8B9300100C13
01798A330F3C5863
014D0A33002A1A13
000A2903FFCA2483
41990AB30044AC83
000C8413001ABA93
0004A40301991663
00042783FFE47413
040790630017F793
008A202300098593
DF5FF0EF000D0513
001989930004A783
00F4A023FFE7F793
000A248300042783
00F420230017E793
07990463012A2223
00042A030044A403
FFEA7A1300442703
000A2783000A0863
140784630017F793
0007278300070863
080788630017F793
0000061301691A63
00048513000A8593
00042783CD9FF0EF
00F42023FFE7F793
0017F7130004A783
FFF9899300070C63
0004A403F29FF06F
F99FF06FFFE47413
00F4A0230017E793
0281240302C12083
0201290302412483
01812A0301C12983
01012B0301412A83
00812C0300C12B83
00012D0300412C83
0000806703010113
FFE7F79300042783
000A07931080006F
000707930B990863
0016F6930007A683
0004A7030A069263
0009859300042683
FFE6F69300177713
00E4202300D76733
000D05130004A703
00E4A02300176713
001767130007A703
0029979300E7A023
FE87AE2300FD07B3
F5691EE3CB1FF0EF
02C1208302812403
01C1298302012903
01012B0301812A03
00812C0300C12B83
00012D0300412C83
00048513000A8593
0241248301412A83
0301011300000613
000A0793BB9FF06F
00070793F79900E3
01991463F4079CE3
00299B9300070A13
017D0BB3FFCB8B93
014BA223008BA023
000D051300198593
00042783C31FF0EF
00F42023FFE7F793
000BA403000A2783
00FA20230017E793
00442783EF990CE3
F11FF06F012BA023
0005086300052503
0045278300058C63
0000806700079463
FE9FF06F00078513
FFE7F79300052783
FD010113FE9FF06F
0291222302812423
0211262301312E23
01412C2303212023
0161282301512A23
0301041301712623
0005A2230005A783
0017F79300050993
0005278300F5A023
0407966300058493
0010079300B9A023
0005A78300F52423
00F5A0230017E793
02C12083FD040113
0241248302812403
01C1298302012903
01412A8301812A03
00C12B8301012B03
0000806703010113
00010A9300852783
0137879300279793
40F10133FF07F793
000A061300010A13
00251793A91FF0EF
FFC92B8300FA0933
00050B130049A783
00048513000B8593
00154593000780E7
000B851300048613
A3DFF0EF0FF5F593
001B0B130004A783
FFE7F79300992023
000B0B9300F4A023
0010081300090793
000A270301784A63
0017E79300072783
FFC7A6030CC0006F
00062703FFC78913
0A071E6300177713
FF878493FF87A583
000706930045A703
0005A68300E61663
04068063FFE6F693
000487930006A503
0205186300157513
FFEB8B930005A703
00E5A023FFE77713
0017671300062703
0006A70300E62023
00E6A02300176713
002B9793F81FF06F
FFC7A78300FA07B3
40E6073300462683
40D787B300173713
00F708630017B793
000A0513000B8593
FFFB8593A19FF0EF
A0DFF0EF000A0513
000727830004A703
00F720230017E793
0007278300092703
00F72023FFE7F793
0167D4630089A783
000A27830169A423
000A811300F9A023
FD010113E61FF06F
0291222302812423
0161282301412C23
0181242301712623
0321202302112623
01512A2301312E23
0301041301912223
00010B9300852783
0027979300050B13
FF07F79301378793
00010A1340F10133
00058493000A0613
00251C138E1FF0EF
FFCC2783018A0C33
0004A90310979263
FFE9791300050993
0044A7830C090463
001007930C078063
0137D46300000513
012C2023FF8C2503
0049278300198713
0007099300271A93
0E079E63015A0AB3
10050263FF8AAC83
0009061300452583
0015B593409585B3
0F949A63851FF0EF
0004A78300092703
0017F793FFE77713
00F4A02300E7E7B3
0017F79300092783
00F9202300F4E7B3
00F922230044A783
FFCC2783FFCAA703
FEEC2E230004A223
0004A683FEFAAE23
FFE6F79300092703
00F7673300177713
0009278300E4A023
FFE7F7930016F693
00F9202300D7E7B3
FFE7F9130004A783
0044A90300091463
0B374C6300100713
0A090463012B2023
0017E79300092783
000B811300F92023
02C12083FD040113
0241248302812403
01C1298302012903
01412A8301812A03
00C12B8301012B03
00412C8300812C03
0000806703010113
0017071300FAA023
EE9FF06F00078913
F11FF06F012B2023
00048613004CA583
412585B3000C8513
F44FF0EF0015B593
000926830004A703
FFE6F69300177793
00F4A02300D7E7B3
FFE7771300092783
00E7E7B30017F793
000B2423EF5FF06F
00299A93F65FF06F
FF8AA503015A0AB3
0017F79302091863
0607946300048613
0000061300452583
0015B593409585B3
000A2783EE0FF0EF
F29FF06F00FB2023
0009061300452583
0015B593409585B3
0004A783EC0FF0EF
000788630017F793
0017F79300092783
0009278300079A63
00F920230017E793
FF2AAE23FBDFF06F
0009859300000613
8A9FF0EF000A0513
00052503FA5FF06F
0005166300058793
0000806700000513
FFF007130085A683
80DFF06F00E69463
002697130005A603
0007250300E60733
FE0514E300452503
00D585330045A583
00050C6300054503
00D7A423FFF68693
00008067FFC72503
0087A68300E7A423
00D05863FFF68713
0006C68300D586B3
00E7A423FE0684E3
00271713F80748E3
0007250300E60733
FF01011300008067
0005851300050793
0006861300060593
000780E700112623
545020EF091020EF
0000806700000513
00812423FF010113
0450051300050413
0091222300112623
000400E700058493
0520051300048593
00040313000400E7
00C1208300812403
0041248300048593
0101011305200513
0005A78300030067
00F5A02300178793
C947A303000067B7
FB01011300030067
03312E2304812423
03512A2303412C23
0411262303612823
0521202304912223
0381242303712623
03A1202303912223
00050A1301B12E23
0006099300058A93
0010041300068B13
0007041300E05463
02000C1300100793
03000C1300FB1463
001009133B9AD4B7
0000071300A00C93
00200D939FF48493
00148B9300A00D13
0934F26300071463
000A85930379D533
0305051300190913
00100713000A00E7
00100793FFFC8C93
03A4D4B30379F9B3
000A8593FCFC96E3
000A00E703098513
4124043300300793
04C1208306FB0A63
0441248304812403
03C1298304012903
03412A8303812A03
02C12B8303012B03
02412C8302812C03
01C12D8302012D03
0000806705010113
F96DEAE3F9944CE3
000C0513000A8593
000A00E700E12623
00C1270300190913
000A8593F79FF06F
000A00E702000513
FE8048E3FFF40413
000067B7F8DFF06F
00008067C8A7AA23
04812423FB010113
0521202304912223
03412C2303312E23
0391222303512A23
01B12E2303A12023
0361282304112623
0381242303712623
0005849300050413
00068D1300060A93
FFF0091300000A13
00000C9300000993
000AC50380000DB7
04C1208304051063
0441248304812403
03C1298304012903
03412A8303812A03
02C12B8303012B03
02412C8302812C03
01C12D8302012D03
0000806705010113
02500693000C9E63
0004859336D50A63
001A8A93000400E7
06400693FA5FF06F
06A6E26310D50E63
02A6EA6303900693
0ED5746303100693
34D50A6302D00693
0CF5006303000793
02E5126302500713
0250051300048593
15C0006F000400E7
1AD50E6305800693
2EE50E6306300713
0250051300048593
00048593000400E7
FD5FF06F000AC503
16D50A6307000693
0690069302A6E063
06C006930AD50263
0680069308D50A63
FC5FF06FF6D506E3
10D5066307500693
0730071302A6EE63
000D2C03FAE518E3
000C0B93004D0B13
26051863000BC503
00F9986300300793
41790BB3418B8BB3
000B0D1327704663
078006930C80006F
07A0069312D50463
00095E63FA9FF06F
FD05091328098863
00200993F00992E3
FE0948E3EFDFF06F
02D9093300A00693
01250933FD090913
001A0A13FE1FF06F
040A1263EDDFF06F
004D0D13000D2603
0004859302065063
00C1202302D00513
00012603000400E7
40C00633FFF90913
0009869300090713
0004051300048593
03C0006FC95FF0EF
FAEA0EE300100713
FF87F713007D0793
0047268300072603
01B6073300870D13
00D7073300C73733
00048593FA0700E3
BF5FF0EF00040513
E59FF06F00000C93
000D2603000A1863
F9DFF06F004D0D13
FEEA08E300100713
FF87F713007D0793
0007260300870D13
FC0710E300472703
FFF7C793800007B7
FB1FF06FF6C7F8E3
0300051300048593
00048593000400E7
000400E707800513
0010099300800913
0B46C26300100693
00012423000D2783
00F12223004D0D13
00000B9301000C13
0100089300012023
0081258300412503
002B1613FFF88B13
C3CFE0EF01112623
0805186300F57513
0300069300012783
00C1288300079863
08F8966300100793
0185151300A68533
4185551300048593
001B8B93000400E7
00300693040B1863
D6D998E300000C93
41770BB300191713
00048593F17054E3
000400E702000513
FEDFF06FFFFB8B93
FF87F693007D0793
00868D130006A783
0046A78300F12223
F55FF06F00F12423
000B089301912023
00900793F59FF06F
F8A7E2E305700693
F7DFF06F03000693
00F12623FFFC0793
0010079301894C63
0004859300F99C63
000400E703000513
FC1FF06F00C12C03
FEF99AE300200793
0200051300048593
00048593FE5FF06F
000400E7001B8B93
00048593D81FF06F
000400E702000513
D85FF06FFFFB8B93
00048593000D2503
000400E7004D0B13
00000A13D75FF06F
00000993FFF00913
C89FF06F00100C93
C81FF06F00300993
C79FF06F00100993
00050613FE010113
0005869300002537
00C105939D450513
0001262300112E23
01C12083BA1FF0EF
0000806702010113
02B12223FC010113
00112E2302410593
02D1262302C12423
02F12A2302E12823
03112E2303012C23
FA5FF0EF00B12623
0401011301C12083
000065B700008067
FF01011300006537
88C5051385858593
0011262301E00613
000055B7FA9FF0EF
0060051346058593
00008067A99FE0EF
3007A7F300800793
0000806710500073
00A7953300100793
0000806730452573
00A7953300100793
0000806730453573
3007B7F300800793
3440507330405073
FF01011300008067
0091222300812423
0011262300006437
0005049300A00793
00F51C63D0040413
00D0059300042503
0047A78300452783
00042503000780E7
004527830FF4F593
000780E70047A783
0081240300C12083
0041248300048513
0000806701010113
0645051300002537
00006537A65FF06F
89850513FF010113
1EC000EF00112623
D0A7A023000067B7
00C12083FD9FF0EF
0101011300000513
FF01011300008067
0011262300700513
800016B7F31FF0EF
0003D7370186A783
00E787B309070713
00F6AC2300700513
00C12083F01FF0EF
0101011300100513
FF0101134450206F
0011262300700513
800016B7EF1FF0EF
0003D7370186A783
00E787B309070713
00F6AC2300700513
00C12083EC1FF0EF
0101011300000513
0000806700008067
0000806700000513
0005C70300054783
0007966300E79463
0000806740E78533
0015859300150513
0FF5F693FE1FF06F
0037F71300050793
0FF5F59304071863
00B765B300859713
00B765B301059713
0007871300C78333
40E308B300300813
0026571303186E63
00B787B300271593
02B70733FFC00593
00E7873300C70733
0000806702E79463
00178793FE060EE3
FFF60613FED78FA3
00470713F9DFF06F
FB9FF06FFEB72E23
FED78FA300178793
800017B7FD1FF06F
0000806700B78423
0087C783800017B7
00F5802300000513
0000051300008067
0025171300008067
00150513000067B7
002515138C078793
00E78733FF010113
0081242300A787B3
0007240300912223
001126230007A483
00C1208300946C63
0041248300812403
0000806701010113
0004051300042783
000780E70047A783
0004222300050463
FCDFF06F00C40413
000067B7FF010113
000064B700912223
0011262300812423
01212023CA878413
CD848493CA878793
0005091300941C63
0294146300078413
0440006F00000413
0007086300442703
0007270300042703
00C4041302A70863
00442783FD1FF06F
00C4041300079663
00042783FCDFF06F
0007A58300090513
FE0514E3E49FF0EF
00C1208300040513
0041248300812403
0101011300012903
FF01011300008067
0011262300812423
300437F300800413
00A04463025020EF
0010059300100513
C8DFF0EF0F1020EF
00006537FE5FF06F
CF050613000067B7
40C7863315078793
CF05051300000593
FF010113DFDFF06F
0011262300200513
00006537E9DFF0EF
BDDFF0EF8D450513
E89FF0EF00300513
D30FE0EF1F8020EF
0AC78793000067B7
FFE7771300C7C703
00C1208300E78623
0000806701010113
08812C23F6010113
00006437000087B7
1507879309312623
00F9A22311C40993
0700061301010793
0007851300000593
08912A2308112E23
D71FF0EF09212823
00A9A42300100713
00E10EA300000513
00100513E0DFF0EF
10100793E05FF0EF
1CD010EF00F11E23
90478793000067B7
00F1222300006937
00100793000026B7
0AC90493000075B7
0000071300F12023
0000089300000793
3BC6869300000813
3505859340000613
0299A0230AC90513
00D4C7835A1010EF
FFB7F71311C40413
01B7F79300E486A3
0184A78300079A63
0AC9051300079663
000067B7134010EF
00F1222390C78793
0010079300006537
000075B7000026B7
00F1202303C50493
0000081302800893
0000071300000793
2000061336C68693
03C5051375058593
00D4C783531010EF
0080051300942623
00F486A3FFB7F793
13478793000067B7
00F42E2300F42C23
0085751330053573
000067B7CD1FD0EF
FF01011311C7A703
0011262300812423
0007841300912223
000064B702070E63
00006537000065B7
10000693A1858593
804505139F448613
00006537A19FF0EF
A0DFF0EFA3050513
9F44851310000593
11C40793A3DFF0EF
00F7C7030087A783
02F71E6300100793
000065B700006437
A345859300006537
9F44061310100693
9CDFF0EF80450513
A305051300006537
101005939C1FF0EF
9F1FF0EF9F440513
11C78793000067B7
00F747830087A703
00F707A3FFF78793
0081240300C12083
0101011300412483
0005242300008067
00A5202300052623
0000806700A52223
02812423FD010113
0005041301412C23
0291222302112623
01312E2303212023
00058A1301512A23
00C42703EF5FF0EF
11C78793000067B7
0084260302070063
04D60E630087A683
609000EF060A1063
0280006FFF000513
00E686830087A683
001707130087A783
00E4262300D42823
5E1000EF00F42423
02C1208300000513
0241248302812403
01C1298302012903
01412A8301812A03
0000806703010113
FBDFF06F01042683
00E6890300E60783
000789130127D463
0000091300095463
3009B9F300800993
D0448513000064B7
411010EF0089F993
00006AB702051E63
00006537000065B7
04E0069393058593
80450513914A8613
00006537879FF0EF
86DFF0EF94850513
914A851304E00593
D044851389DFF0EF
00842503425010EF
00F9566300E50783
558010EF00090593
00040613000A0693
D044851300098593
00A126234BC010EF
509000EF00051863
F29FF06F00C12503
0104298300042783
00078C6300F40E63
0137D46300E78783
0009D46300078993
0080091300000993
D044851330093973
359010EF00897913
00006A3702051E63
00006537000065B7
04E0069393058593
80450513914A0613
00006537FC0FF0EF
FB4FF0EF94850513
914A051304E00593
D0448513FE4FF0EF
0084250336D010EF
00F9866300E50783
4A0010EF00098593
321010EFD0448513
0000643702051E63
00006537000065B7
0610069396058593
8045051391440613
00006537F60FF0EF
F54FF0EF97850513
9144051306100593
30092973F84FF0EF
FF500513425000EF
00C52783E45FF06F
00812C23FE010113
00912A2300112E23
0131262301212823
02079E6300050413
000065B7000064B7
9BC5859300006537
98C486130D400693
EF4FF0EF80450513
A305051300006537
0D400593EE8FF0EF
F18FF0EF98C48513
00842703000067B7
02F70E631247A783
000065B7000064B7
9D45859300006537
98C486130D500693
EACFF0EF80450513
A305051300006537
0D500593EA0FF0EF
ED0FF0EF98C48513
00C42783C3DFF0EF
02E7846300100713
00F42623FFF78793
01C1208301812403
0101290301412483
0201011300C12983
008004933450006F
000069373004B4F3
0084F493D0490513
02051E631BD010EF
000065B7000069B7
9305859300006537
9149861304E00693
E24FF0EF80450513
9485051300006537
04E00593E18FF0EF
E48FF0EF91498513
1D1010EFD0490513
0104258300842503
00F5846300E50783
00040513304010EF
00A424236C0000EF
06050A6300050993
01F7F79300D54783
0185278300079863
429000EF00079463
159010EFD0490513
0000693702051E63
00006537000065B7
0610069396058593
8045051391490613
00006537D98FF0EF
D8CFF0EF97850513
9149051306100593
3004A4F3DBCFF0EF
0609A62300E98783
EF5FF06F00F42823
D049051300042623
02051E630FD010EF
000065B700006437
9605859300006537
9144061306100693
D3CFF0EF80450513
9785051300006537
06100593D30FF0EF
D60FF0EF91440513
EA5FF06F3004A4F3
01F7F79300D54783
0185250300079863
0000806700153513
0000806700000513
00E5868300E50703
00D74C6300100793
00E6C86300000793
0105A50301052783
0007851300A7B7B3
FF01011300008067
E9CFF0EF00112623
D107A783000067B7
0000673700C12083
12A7262300A78533
0007851300000593
16C0206F01010113
FF01011300052783
0011262300812423
0005041300912223
000064B702079863
00006537000065B7
80450513AB458593
A844861318300693
18300593C60FF0EF
C90FF0EFA8448513
00C1208300042503
0041248300812403
0000806701010113
00812C23FE010113
0141242301212823
00912A2300112E23
0005091301312623
0080041300058A13
000064B730043473
00847413D0848513
02051E63774010EF
000065B7000069B7
9305859300006537
9149861304E00693
BDCFF0EF80450513
9485051300006537
04E00593BD0FF0EF
C00FF0EF91498513
788010EFD0848513
1207A623000067B7
00A0079300990913
000067B702F94933
000067B7D127A823
EC9FF0EFD147A623
728010EFD0848513
000064B702051E63
00006537000065B7
0610069396058593
8045051391448613
00006537B68FF0EF
B5CFF0EF97850513
9144851306100593
30042473B8CFF0EF
0181240301C12083
0101290301412483
00812A0300C12983
0000806702010113
00812C23FE010113
00112E2301212823
0131262300912A23
0080041300050913
000064B730043473
00847413D0848513
02051E6366C010EF
000065B7000069B7
9305859300006537
9149861304E00693
AD4FF0EF80450513
9485051300006537
04E00593AC8FF0EF
AF8FF0EF91498513
680010EFD0848513
E15FF0EF00890513
2F0000EF00090593
D084851300D94783
00F906A3FFD7F793
02051E6362C010EF
000065B7000064B7
9605859300006537
9144861306100693
A6CFF0EF80450513
9785051300006537
06100593A60FF0EF
A90FF0EF91448513
01C1208330042473
0009242301812403
0101290301412483
0201011300C12983
000067B700008067
FF01011311C7A783
0011262300812423
0005841300912223
5A8010EF04079E63
000064B702051E63
00006537000065B7
0780069396058593
8045051391448613
000065379E8FF0EF
9DCFF0EF97850513
9144851307800593
00040513A0CFF0EF
00C1208300812403
0101011300412483
550010EFC30FD06F
000064B702051E63
00006537000065B7
0610069396058593
8045051391448613
00006537990FF0EF
984FF0EF97850513
9144851306100593
008474139B4FF0EF
00C1208330042473
0041248300812403
0000806701010113
11C7270300006737
BC4FD06F00071463
3007A7F300857793
0080051300008067
0085751330053573
FE010113FD9FF06F
00112E2300812C23
0121282300912A23
0080041301312623
000064B730043473
00847413D0848513
02051E63474010EF
000065B700006937
9305859300006537
9149061304E00693
8DCFF0EF80450513
9485051300006537
04E005938D0FF0EF
900FF0EF91490513
00006937D0848513
11C92783484010EF
02078E6311C90913
000065B7000069B7
A185859300006537
9F49861310000693
88CFF0EF80450513
A305051300006537
10000593880FF0EF
8B0FF0EF9F498513
00F7C70300892783
02F71E6300100793
000065B7000069B7
A345859300006537
9F49861310100693
844FF0EF80450513
A305051300006537
10100593838FF0EF
868FF0EF9F498513
00F7478300892703
00F707A3FFF78793
3B0010EFD0848513
000064B702051E63
00006537000065B7
0610069396058593
8045051391448613
00006537FF1FE0EF
FE5FE0EF97850513
9144851306100593
30042473814FF0EF
0181240301C12083
0101290301412483
0201011300C12983
000067B700008067
FF010113CA47A783
0011262300812423
0005841300912223
000064B702F59863
00006537000065B7
80450513B3858593
A844861328C00693
28C00593F79FE0EF
FA9FE0EFA8448513
0004278300442703
0041248300C12083
00E7A22300F72023
0004222300042023
0101011300812403
0005278300008067
0000079300F51463
0000806700078513
01212823FE010113
00112E2301312623
00912A2300812C23
0080091300050993
000064B730093973
00897913D0848513
02051E6326C010EF
000065B700006437
9305859300006537
9144061304E00693
ED5FE0EF80450513
9485051300006537
04E00593EC9FE0EF
EF9FE0EF91440513
280010EFD0848513
F71FF0EF00098513
D084851300050413
02051E6323C010EF
000065B7000069B7
9605859300006537
9149861306100693
E7DFE0EF80450513
9785051300006537
06100593E71FE0EF
EA1FE0EF91498513
0C04066330092973
3009397300800913
00897913D0848513
02051E631BC010EF
000065B7000069B7
9305859300006537
9149861304E00693
E25FE0EF80450513
9485051300006537
04E00593E19FE0EF
E49FE0EF91498513
1D0010EFD0848513
965FF0EF00840513
E41FF0EF00040593
D084851300D44783
00F406A3FFD7F793
02051E6317C010EF
000065B7000064B7
9605859300006537
9144861306100693
DBDFE0EF80450513
9785051300006537
06100593DB1FE0EF
DE1FE0EF91448513
0004242330092973
091010EF01840513
01C1208300040513
0141248301812403
00C1298301012903
0000806702010113
02812423FD010113
0321202302912223
01312E2302112623
000067B703010413
00050493CA47A783
02F5986300058913
000065B7000069B7
B385859300006537
2B00069380450513
D25FE0EFA8498613
A84985132B000593
00C4A703D55FE0EF
00F4A62300170793
04079A6300E92823
002797130084A783
FF07771301770713
40E1013301778793
00F10713FF07F793
00F1079340F10133
FF077713FF07F793
FFF00793FCF42C23
FCF42E23FCE42A23
00048513FD440593
02051863DD4FE0EF
0004851300090593
FD04011391CFE0EF
0281240302C12083
0201290302412483
0301011301C12983
00C4A78300008067
00E4A62300178713
FB5FF06F00F52823
CA47A783000067B7
00812423FF010113
0011262300912223
0005041301212023
02F5986300058493
000065B700006937
B385859300006537
2CB0069380450513
C2DFE0EFA8490613
A84905132CB00593
00048593C5DFE0EF
A90FE0EF00040513
0007946300042783
00C1208300042623
0041248300812403
0101011300012903
0000059300008067
FF010113830FE06F
0000643700812423
0005091301212023
0245051311C40513
0011262300912223
11C40413FD5FF0EF
0005146300050493
06091E6300C42483
02079E6300842783
000065B700006937
ACC5859300006537
A849061307F00693
B85FE0EF80450513
A305051300006537
07F00593B79FE0EF
BA9FE0EFA8490513
00D7C70300842783
0207166301F77713
07F0071300E7D683
02F4202302D77063
0081240300C12083
0001290300412483
0000806701010113
0097846300842783
02942023E5CFF0EF
FE010113FD9FF06F
0000693701212823
0087A78311C90793
00812C2300112E23
00912A2300F7C783
11C9091301312623
0000643702079E63
00006537000065B7
22100693A5C58593
80450513A8440613
00006537AD1FE0EF
AC5FE0EFA3050513
A844051322100593
00092783AF5FE0EF
0000643702078E63
00006537000065B7
22200693A1858593
80450513A8440613
00006537A91FE0EF
A85FE0EFA3050513
A844051322200593
00800413AB5FE0EF
000064B730043473
00847413D0848513
02051E635D5000EF
000065B7000069B7
9305859300006537
9149861304E00693
A3DFE0EF80450513
9485051300006537
04E00593A31FE0EF
A61FE0EF91498513
5E9000EFD0848513
0010051300892703
0017879300F74783
E21FF0EF00F707A3
599000EFD0848513
000064B702051E63
00006537000065B7
0610069396058593
8045051391448613
000065379D9FE0EF
9CDFE0EF97850513
9144851306100593
300424739FDFE0EF
01C1208301812403
0101290301412483
0201011300C12983
FE010113865FF06F
0121282300812C23
00912A2300112E23
0005091301312623
3004347300800413
D0848513000064B7
4E1000EF00847413
000069B702051E63
00006537000065B7
04E0069393058593
8045051391498613
00006537949FE0EF
93DFE0EF94850513
9149851304E00593
D084851396DFE0EF
000065374F5000EF
1405051300090593
00D94783BA9FF0EF
0407E79300000513
D21FF0EF00F906A3
499000EFD0848513
000064B702051E63
00006537000065B7
0610069396058593
8045051391448613
000065378D9FE0EF
8CDFE0EF97850513
9144851306100593
300424738FDFE0EF
0181240301C12083
0101290301412483
0201011300C12983
FF05278300008067
00812C23FE010113
00112E2301312623
0121282300912A23
0005041301412423
0C078463FE850993
3004B4F300800493
D089051300006937
3D1000EF0084F493
00006A3702051E63
00006537000065B7
04E0069393058593
80450513914A0613
00006537839FE0EF
82DFE0EF94850513
914A051304E00593
D089051385DFE0EF
FF0405133E5000EF
00098593B78FF0EF
FF544783855FF0EF
FFD7F793D0890513
391000EFFEF40AA3
0000693702051E63
00006537000065B7
0610069396058593
8045051391490613
00006537FD0FE0EF
FC4FE0EF97850513
9149051306100593
3004A4F3FF4FE0EF
FF544783FE042823
FEB7F79300098513
A84FF0EFFEF40AA3
0181240302050463
0141248301C12083
00812A0301012903
00C1298300098513
DD9FF06F02010113
0181240301C12083
0101290301412483
00812A0300C12983
0000806702010113
00812C23FE010113
00112E2301312623
0121282300912A23
0005099301412423
3004347300800413
D0848513000064B7
291000EF00847413
0000693702051E63
00006537000065B7
04E0069393058593
8045051391490613
00006537EF8FE0EF
EECFE0EF94850513
9149051304E00593
00006937F1CFE0EF
11C90913D0848513
02490A1329D000EF
000A051300098593
00098593A51FF0EF
945FF0EF000A0513
0089250300D9C783
413505330407E793
00F986A300153513
D0848513AB5FF0EF
02051E6322D000EF
000065B7000064B7
9605859300006537
9144861306100693
E6CFE0EF80450513
9785051300006537
06100593E60FE0EF
E90FE0EF91448513
01C1208330042473
0141248301812403
00C1298301012903
0201011300812A03
000067B700008067
06078663D107A783
11C78793000067B7
07F006930087A703
04C6EA6300E75603
00E70603000066B7
04D64263D0C6A683
CA46A683000066B7
0187268302D70C63
0107A68302069863
FF01011302D54063
0011262300070513
00C12083E81FF0EF
8F8FF06F01010113
00D7A82340A686B3
FE01011300008067
0131262300812C23
00912A2300112E23
0005099301212823
3004347300800413
D0848513000064B7
0F9000EF00847413
0000693702051E63
00006537000065B7
04E0069393058593
8045051391490613
00006537D60FE0EF
D54FE0EF94850513
9149051304E00593
D0848513D84FE0EF
00D9C78310D000EF
11C9091300006937
00078E630407F793
0249051300098593
00D9C7838B1FF0EF
00F986A3FBF7F793
4135053300892503
921FF0EF00153513
099000EFD0848513
000064B702051E63
00006537000065B7
0610069396058593
8045051391448613
00006537CD8FE0EF
CCCFE0EF97850513
9144851306100593
30042473CFCFE0EF
0181240301C12083
0101290301412483
0201011300C12983
FE01011300008067
00912A2300812C23
0121282300050413
0131262300112E23
0006091300058493
00D44783EC5FF0EF
00F406A30027E793
000067B706048663
00942423CA47A783
000069B702F41863
00006537000065B7
80450513B3858593
A849861327600693
27600593C38FE0EF
C68FE0EFA8498513
06F48C630004A783
00E4070306078A63
04D75C6300E78683
00F420230047A703
0087202300E42223
FFF007930087A223
0099091306F90463
02C9463300A00613
0181240301840513
0141248301C12083
00C1298301012903
71458593000035B7
0016061302010113
0044A6834910006F
0007A78300D78663
0044A783F8079CE3
00F4222300942023
0087A0230044A783
F99FF06F0084A223
0181240301C12083
0101290301412483
0201011300C12983
FF01011300008067
00812423000067B7
1247A50300050413
0005849300912223
0006861300060593
EB1FF0EF00112623
6E0000EF00040513
0000643702051E63
00006537000065B7
0780069396058593
8045051391440613
00006537B20FE0EF
B14FE0EF97850513
9144051307800593
00812403B44FE0EF
0004851300C12083
0101011300412483
FE010113D68FC06F
0121282300812C23
00112E2301312623
0141242300912A23
0005091301512223
0080041300058993
000064B730043473
00847413D0848513
02051E63624000EF
000065B700006A37
9305859300006537
914A061304E00693
A8CFE0EF80450513
9485051300006537
04E00593A80FE0EF
AB0FE0EF914A0513
638000EFD0848513
D4DFE0EF00090513
00050A9301899993
0A0508634189D993
140A0A1300006A37
000A051300090593
000A0513DD0FF0EF
0009059301390723
00100513CC0FF0EF
D0848513E44FF0EF
02051E635BC000EF
000065B7000064B7
9605859300006537
9144861306100693
9FCFE0EF80450513
9785051300006537
061005939F0FE0EF
A20FE0EF91448513
040A806330042473
1247A783000067B7
0207986300F7C783
01C1208301812403
0101290301412483
00812A0300C12983
0201011300412A83
0139072386CFF06F
01C12083F7DFF06F
0141248301812403
00C1298301012903
00412A8300812A03
0000806702010113
00003737000067B7
AB87071311C78793
0000051300000593
0207A6230207A223
02E7A4230207A823
00E50503D19FE06F
FE01011300008067
0000643700812C23
00112E2311C42783
0121282300912A23
11C4041301312623
000064B702078E63
00006537000065B7
37E00693A1858593
80450513A8448613
00006537900FE0EF
8F4FE0EFA3050513
A844851337E00593
000067B7924FE0EF
CA47A78300842703
008007930CF70663
000064B73007B7F3
0087F993D0848513
02051E63434000EF
000065B700006937
9305859300006537
9149061304E00693
89CFE0EF80450513
9485051300006537
04E00593890FE0EF
8C0FE0EF91490513
448000EFD0848513
0244091300842583
BFCFF0EF00090513
0009051300842583
00100513AF0FF0EF
D0848513C74FF0EF
02051E633EC000EF
000065B700006437
9605859300006537
9144061306100693
82CFE0EF80450513
9785051300006537
06100593820FE0EF
850FE0EF91440513
008005133009A7F3
0181240330053573
0141248301C12083
00C1298301012903
0201011300857513
FD010113A60FC06F
000064B702912223
0281242311C4A783
0321202302112623
01412C2301312E23
11C4849300050413
0000693702078E63
00006537000065B7
39900693A1858593
80450513A8490613
00006537F99FD0EF
F8DFD0EFA3050513
A849051339900593
FFF00793FBDFD0EF
000069371AF41263
00006537000065B7
39A00693AEC58593
80450513A8490613
00006537F59FD0EF
F4DFD0EFA3050513
A849051339A00593
00A00793F7DFD0EF
02F4443300940413
00800993765000EF
0014041300012623
3009B9F300A40933
0089F99300C10513
02051E63284000EF
000065B700006A37
9305859300006537
914A061304E00693
EEDFD0EF80450513
9485051300006537
04E00593EE1FD0EF
F11FD0EF914A0513
298000EF00C10513
911FF0EF0084A503
000035B70084A503
0185051300040613
77C000EF71458593
00C105130084A703
0107E79300D74783
230000EF00F706A3
0000643702051E63
00006537000065B7
0780069396058593
8045051391440613
00006537E71FD0EF
E65FD0EF97850513
9144051307800593
00098513E95FD0EF
0084A7838C8FC0EF
0107F79300D7C783
0000643702078E63
00006537000065B7
3B700693B0058593
80450513A8440613
00006537E21FD0EF
E15FD0EFA3050513
A84405133B700593
639000EFE45FD0EF
0000041340A90533
3E80079302A05663
0640061302F515B3
02F5053300000693
000504138E0FC0EF
E8041CE300C0006F
00040513C8DFF0EF
0281240302C12083
0201290302412483
01812A0301C12983
0000806703010113
1247A503000067B7
00D5478300008067
0007986301F7F793
0015351301852503
0000051300008067
000067B700008067
00A0353311C7A503
000067B700008067
00C7C5031247A783
0000806700157513
02012303FE010113
00112E2300812C23
0005041300612023
000067B7A35FC0EF
01C120831247A783
06F424230687A783
0201011301812403
0605278300008067
00812423FF010113
0005041300112623
000780E700078463
F61FF0EF00040513
0004051302050463
00D44783F3CFF0EF
0087E79300C12083
0081240300F406A3
0000806701010113
0027F79300D44783
0004051300078663
01842783999FE0EF
01840513FC0786E3
FC1FF06F7AC000EF
00C506A300D50623
000507A300B50723
00052E2300052C23
0005250300008067
000067B700050E63
003575131307C783
00A0353340F50533
0010051300008067
000067B700008067
0147C70311C78793
00E7E7B30087A783
00F7186300052703
0010051300052023
0000051300008067
000067B700008067
0147C70311C78793
00E7E7B30087A783
0000806700F52023
00812C23FE010113
00112E2301212823
0131262300912A23
0080041300050913
000064B730043473
00847413D1448513
02051E63F5DFF0EF
000065B7000069B7
9305859300006537
9149861304E00693
BC5FD0EF80450513
9485051300006537
04E00593BB9FD0EF
BE9FD0EF91498513
F71FF0EFD1448513
0047F71300D94783
D144851306071463
02051E63F2DFF0EF
000065B7000064B7
9605859300006537
9144861306100693
B6DFD0EF80450513
9785051300006537
06100593B61FD0EF
B91FD0EF91448513
01C1208330042473
0141248301812403
00C1298301012903
0000806702010113
00F906A3FFB7F793
D89FF0EF00090513
0009051300050663
0004059397CFF0EF
01C1208301812403
00C1298301012903
01412483D1448513
8C9FE06F02010113
03512223FC010113
000066B700068A93
02812C2311C6A683
0331262302912A23
02112E2303412423
0005049303212823
00060A1300058993
04068E6304412403
000065B700006937
1B20069300006537
A1858593B4C90613
01112E2380450513
00F12A2301012C23
A85FD0EF00E12823
B805051300006537
1B200593A79FD0EF
AA9FD0EFB4C90513
0181280301C12883
0101270301412783
0001222304012683
00D12023000A0613
000A869300098593
CE5FF0EF00048513
00F40863FFF00793
0004851302041A63
03C12083E11FF0EF
0004851303812403
0341248303012903
02812A0302C12983
0401011302412A83
0094041300008067
02C4463300A00613
71458593000035B7
0016061301848513
FB9FF06F2B0000EF
000067B7FD010113
0000693703212023
0291222302812423
01312E2302112623
CD87841301412C23
CD890913CD878493
0004841303246E63
FFF00493875FE0EF
00003A3700A00993
0281240307246463
0241248302C12083
01C1298302012903
0301011301812A03
02C42783E55FE06F
0204278300F12223
0144278300F12023
0184280301C42883
00C4268301042703
0044258300842603
BE5FF0EF00042503
0487AE2300042783
F85FF06F03040413
0096086302442603
0006186300042503
03040413D01FF0EF
00960613F81FF06F
714A059303364633
0016061301850513
FE1FF06F1C8000EF
00812C23FE010113
00112E2300912A23
0005049301212823
0080041300012623
00C1051330043473
C39FF0EF00847413
0000693702051E63
00006537000065B7
04E0069393058593
8045051391490613
000065378A1FD0EF
895FD0EF94850513
9149051304E00593
00C105138C5FD0EF
00C4C783C4DFF0EF
02078E630017F793
000065B700006937
BE05859300006537
BA89061302900693
855FD0EF80450513
C145051300006537
02900593849FD0EF
879FD0EFBA890513
B19FF0EF00048513
00C1051300040593
01C12083DFCFE0EF
0141248301812403
0201011301012903
000067B700008067
00079463D187A783
000005139D9FD06F
0005278300008067
0000673702050263
00E50C63C9C72703
0087A70300078A63
00D7073300852683
0045270300E7A423
00E7A22300F72023
0005222300052023
000067B700008067
FF010113D207C783
0081242300112623
FFF0051300912223
8000053700079663
000067B7FFF54513
0007A403C9878793
0204026302F40463
F69FF0EF00842483
0000051340A484B3
008424030004C863
40A40533F55FF0EF
12C7A783000067B7
00A7D46300078663
00C1208300078513
0041248300812403
0000806701010113
FD01011300052783
0291222302812423
0211262301312E23
01412C2303212023
0161282301512A23
0181242301712623
0005899300050413
02078E6300060493
000065B700006937
C645859300006537
C309061304D00693
ED4FD0EF80450513
A305051300006537
04D00593EC8FD0EF
EF8FD0EFC3090513
0090446301342623
0080099300100493
00006A373009B9F3
0089F993D1CA0513
02051E63A0DFF0EF
000065B700006937
9305859300006537
9149061304E00693
E74FD0EF80450513
9485051300006537
04E00593E68FD0EF
E98FD0EF91490513
A21FF0EFD1CA0513
00950533E45FF0EF
C984A903000064B7
C984849300A42423
00006AB700990C63
00006BB700006B37
0209106300006C37
009420230044A783
0044A78300F42223
0084A2230087A023
0089278305C0006F
C84B05930207D663
C30A861305600693
DECFD0EF804B8513
DE4FD0EFA30C0513
C30A851305600593
00892703E14FD0EF
0AE7D86300842783
00F9242340F707B3
0124202300492783
0087A02300F42223
0004A78300892223
00F4186300978A63
00000593DEDFF0EF
D1CA0513F6CFD0EF
02051E6392DFF0EF
000065B700006437
9605859300006537
9144061306100693
D6CFD0EF80450513
9785051300006537
06100593D60FD0EF
D90FD0EF91440513
02C120833009A9F3
0241248302812403
01C1298302012903
01412A8301812A03
00C12B8301012B03
0301011300812C03
40E787B300008067
0044A78300F42423
00092903EF2788E3
FE010113EE5FF06F
0131262300812C23
00912A2300112E23
0005099301212823
3004347300800413
D1C48513000064B7
849FF0EF00847413
0000693702051E63
00006537000065B7
04E0069393058593
8045051391490613
00006537CB0FD0EF
CA4FD0EF94850513
9149051304E00593
D1C48513CD4FD0EF
0009A78385DFF0EF
00078863FEA00913
C89FF0EF00098513
D1C4851300000913
02051E6380DFF0EF
000065B7000064B7
9605859300006537
9144861306100693
C4CFD0EF80450513
9785051300006537
06100593C40FD0EF
C70FD0EF91448513
01C1208330042473
0009051301812403
0101290301412483
0201011300C12983
FF01011300008067
0011262300812423
0121202300912223
3004347300800413
D1C48513000064B7
F58FF0EF00847413
0000693702051E63
00006537000065B7
04E0069393058593
8045051391490613
00006537BC0FD0EF
BB4FD0EF94850513
9149051304E00593
D1C48513BE4FD0EF
BE9FF0EFF6CFF0EF
D1C4851300050913
02051E63F2CFF0EF
000065B7000064B7
9605859300006537
9144861306100693
B6CFD0EF80450513
9785051300006537
06100593B60FD0EF
B90FD0EF91448513
00C1208330042473
0009051300812403
0001290300412483
0000806701010113
00812C23FE010113
0141242301212823
00912A2300112E23
0005091301312623
0080041300058A13
000064B730043473
00847413D1C48513
02051E63E6CFF0EF
000065B7000069B7
9305859300006537
9149861304E00693
AD4FD0EF80450513
9485051300006537
04E00593AC8FD0EF
AF8FD0EF91498513
E80FF0EFD1C48513
00A95C63AFDFF0EF
00A7D86300100793
00090513000A0593
D1C48513C6CFD0EF
02051E63E2CFF0EF
000065B7000064B7
9605859300006537
9144861306100693
A6CFD0EF80450513
9785051300006537
06100593A60FD0EF
A90FD0EF91448513
01C1208330042473
0141248301812403
00C1298301012903
0201011300812A03
FD01011300008067
01412C2302812423
0291222302112623
01312E2303212023
0161282301512A23
0181242301712623
01A1202301912223
0080041300050A13
30043473BC5FE0EF
D1C9051300006937
D50FF0EF00847413
000064B702051E63
00006537000065B7
04E0069393058593
8045051391448613
000065379B8FD0EF
9ACFD0EF94850513
9144851304E00593
000069B79DCFD0EF
D60FF0EFD1C90513
D149AC23000064B7
D189899300006A37
CF048493C98A0A13
00006BB700006AB7
00006C3700006B37
000A2D0300006CB7
0004A6830009A783
014D0C630044A503
008D2703000D0A63
40F707330AE7DC63
00D786B300ED2423
00A7073341F7D713
00E787B300F6B7B3
00F4A22300D4A023
969FF0EF0009A023
AE8FD0EF00000593
CA8FF0EFD1C90513
000064B702051E63
00006537000065B7
0610069396058593
8045051391448613
000065378E8FD0EF
8DCFD0EF97850513
9144851306100593
3004247390CFD0EF
0281240302C12083
0201290302412483
01812A0301C12983
01012B0301412A83
00812C0300C12B83
00012D0300412C83
0000806703010113
41F7559300D706B3
00E6B63300A585B3
40E787B300B60633
000D2423000D0513
00C4A22300D4A023
871FF0EF00F9A023
BF8FF0EFD1C90513
960B859302051663
914A861306100693
844FD0EF804B0513
83CFD0EF978C0513
914A851306100593
3004247386CFD0EF
000D051300CD2783
000780E700800413
D1C9051330043473
B80FF0EF00847413
930C859302051863
914A861304E00693
FF5FC0EF804B0513
9485051300006537
04E00593FE9FC0EF
818FD0EF914A8513
BA0FF0EFD1C90513
000067B7E6DFF06F
00008067CF07A503
CF07A783000067B7
FF0101133E800513
0640061302F535B3
0011262300000693
A9CFB0EF02F50533
0101011300C12083
FF01011300008067
0091222300812423
000064B700006437
CD84041300112623
00946E63CD848493
0081240300C12083
0000051300412483
0000806701010113
0004051301440793
00F42C2300F42A23
01C40413DD9FB0EF
00008067FCDFF06F
00000C1C00000000
00000C1C00000000
00000C1C00000000
00000C1C00000000
00000C1C00000000
00000C1C00000000
00000C1C00000000
0000210400000000
000020D40000545C
000058A000000000
0000000000002144
0000225C00005898
0000545C00000000
0000000000005024
0303030302020100
0404040404040404
0505050505050505
0505050505050505
0606060606060606
0606060606060606
0606060606060606
0606060606060606
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
00005D3800005D24
00005D6000005D4C
00005D8800005D74
007365786574756D
0063696D616E7964
35315B1B4A325B1B
206F6D654448313B
7470697263736544
2D2D2D2D0A6E6F69
2D2D2D2D2D2D2D2D
206E410A2D2D2D2D
6E656D656C706D69
6F206E6F69746174
756C6F7320612066
206F74206E6F6974
696E694420656874
6F6C69685020676E
0A73726568706F73
206D656C626F7270
7373616C63206128
69746C756D206369
206461657268742D
6E6F7268636E7973
206E6F6974617A69
296D656C626F7270
7020736968540A2E
616C756369747261
6D656C706D692072
6E6F697461746E65
74736E6F6D656420
6874207365746172
2065676173752065
69746C756D20666F
656572700A656C70
20656C626974706D
706F6F6320646E61
2065766974617265
2073646165726874
656666696420666F
69727020676E6972
2C7365697469726F
6C6C65770A736120
2520732520736120
687420646E612073
656C732064616572
000A2E676E697065
5320202020202020
20474E4956524154
0000202020202020
49444C4F48202020
4620454E4F20474E
00002020204B524F
474E495441452020
64257325205B2020
0000205D20736D20
50504F5244202020
4620454E4F204445
00002020204B524F
4E494B4E49485420
64257325205B2047
0000205D20736D20
0000005000000043
4864253B64255B1B
6C69685000000000
20726568706F736F
253A73255B206425
000000205D642573
00000BAC00000AF4
00000AE800000BAC
00000B9400000AF4
000054B000000BA0
000054EC000054D0
0000550C00005500
6E6B6E7500005524
65637845006E776F
6163206E6F697470
2820732520657375
000000000A296425
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
7463757274736E49
72646461206E6F69
6173696D20737365
000064656E67696C
7463757274736E49
65636341206E6F69
746C756166207373
656C6C4900000000
74736E69206C6167
006E6F6974637572
696F706B61657242
64616F4C0000746E
7373657264646120
67696C6173696D20
64616F4C0064656E
2073736563636120
000000746C756166
72654B202A2A2A2A
6F6C6C41206C656E
46206E6F69746163
20216572756C6961
0000000A2A2A2A2A
654B202A2A2A2A2A
504F4F206C656E72
2A2A2A2A2A202153
2A2A2A2A0000000A
6C656E72654B202A
202163696E615020
00000A2A2A2A2A2A
6B6E55202A2A2A2A
746146206E776F6E
726F727245206C61
2A2A2A2021642520
7272754300000A2A
6572687420746E65
203D204449206461
746C7561460A7025
74736E6920676E69
206E6F6974637572
2073736572646461
200A78257830203D
257830203A617220
30203A7067202078
3A70742020782578
7420207825783020
0A78257830203A30
7830203A31742020
203A327420207825
3374202078257830
202078257830203A
78257830203A3474
30203A357420200A
3A36742020782578
6120207825783020
2078257830203A30
257830203A316120
203A326120200A78
3361202078257830
202078257830203A
78257830203A3461
7830203A35612020
3A366120200A7825
6120207825783020
0A78257830203A37
0052534900000000
6169746E65737365
646165726874206C
6174614600000000
20746C756166206C
5320217325206E69
2E676E696E6E6970
61746146000A2E2E
20746C756166206C
6165726874206E69
6241202170252064
0A2E676E6974726F
7275705300000000
746E692073756F69
6420747075727265
2164657463657465
6425203A51524920
6D6F682F0000000A
702F666F6C6F2F65
2F737463656A6F72
657A2F7672657773
6372612F72796870
3376637369722F68
742F65726F632F32
00632E6461657268
6F69727028282828
3D20292979746972
202626203034203D
6C64695F73695F7A
6461657268745F65
6461657268742828
292929636E75665F
34282828207C7C20
3E202931202D2030
2939322D2828203D
2828202626202929
797469726F697270
2828203D3E202929
262620292939322D
726F697270282820
3D3C202929797469
31202D2030342820
4553534100292929
4146204E4F495452
205D73255B204C49
0A64253A73252040
766E690900000000
6972702064696C61
252820797469726F
6F6C6C61203B2964
676E617220646577
6F74206425203A65
000000000A642520
6C6F2F656D6F682F
656A6F72702F666F
726577732F737463
72796870657A2F76
2F736F2F62696C2F
632E747265737361
7325204000000000
0000000A3A64253A
0000003074726175
636F6C635F737973
000022480000006B
000000000000223C
0000000000000000
00005CCC00005CA8
00005CD800005CD8
2A2A2A2A00005CD8
6E69746F6F42202A
72796870655A2067
6870657A20534F20
34312E31762D7279
2A2A2A2A2A20302E
6E69616D0000000A
656C646900000000
2E2F2E2E00000000
636E692F2E2E2F2E
6970732F6564756C
00682E6B636F6C6E
6C5F6E6970735F7A
696C61765F6B636F
00000000296C2864
6973727563655209
6C6E697073206576
000000000A6B636F
755F6E6970735F7A
61765F6B636F6C6E
0000296C2864696C
20796D20746F4E09
6B636F6C6E697073
6D6F682F00000A21
702F666F6C6F2F65
2F737463656A6F72
657A2F7672657773
72656B2F72796870
6574756D2F6C656E
6574756D00632E78
5F6B636F6C3E2D78
203E20746E756F63
6574756D00005530
72656E776F3E2D78
72656B5F203D3D20
727275632E6C656E
2E2F2E2E00746E65
72656B2F2E2E2F2E
6C636E692F6C656E
6863736B2F656475
00000000682E6465
656E72656B5F2821
64657473656E2E6C
00295530203D2120
72656B5F00000A09
727275632E6C656E
7361623E2D746E65
5F64656863732E65
212064656B636F6C
72656B5F0031203D
727275632E6C656E
7361623E2D746E65
5F64656863732E65
212064656B636F6C
6D6F682F0030203D
702F666F6C6F2F65
2F737463656A6F72
657A2F7672657773
72656B2F72796870
656863732F6C656E
6572687400632E64
657361623E2D6461
5F6465646E65702E
72656B5F00006E6F
727275632E6C656E
28203D2120746E65
292A2064696F7628
6172756400002930
203D21206E6F6974
0000000029312D28
68745F73695F7A21
6174735F64616572
5F287465735F6574
632E6C656E72656B
202C746E65727275
3C3C204C55312828
0029292929342820
656C64695F736921
2964616572687428
6D6F682F00000000
702F666F6C6F2F65
2F737463656A6F72
657A2F7672657773
72656B2F72796870
657268742F6C656E
00000000632E6461
7364616572685409
746F6E2079616D20
6165726320656220
49206E6920646574
000000000A735253
6C6F2F656D6F682F
656A6F72702F666F
726577732F737463
72796870657A2F76
2F6C656E72656B2F
615F646165726874
0000632E74726F62
2D64616572687428
73752E657361623E
6F6974706F5F7265
312828202620736E
3028203C3C204C55
203D3D2029292929
7373650900005530
74206C6169746E65
6261206461657268
00000A646574726F
6C6F2F656D6F682F
656A6F72702F666F
726577732F737463
72796870657A2F76
2F6C656E72656B2F
2E74756F656D6974
7379732100000063
695F65646F6E645F
64656B6E696C5F73
6F6E3E2D6F742628
643E2D7400296564
3D3E20736B636974
0000198000003020
00005C9800005C98
0000603CFFFFFFF5
00000000000050E4
000050D800000000
00000000000058AC
00000000000050C0
000050CC00000000
0000000000000000
00005CD800005CD8
0000000000000000
0000000000000028
