800015B780002537
08000E1301058593
01B00E9301C50623
00300E1301D50023
08700E1301C50623
0005022301C50423
001FFF9301450F83
00054283000F8E63
020FFF9301450F83
00128293FE0F8CE3
0005D30300550023
0065912300130313
800015B7FD1FF06F
0005A02300958593
0000000000000000
