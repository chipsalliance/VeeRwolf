08000E1380002537
01B00E9301C50623
00300E1301D50023
08700E1301C50623
0005022301C50423
03C5859300000597
01C000EF00058283
0005828300158593
0000006FFE029AE3
00958593800015B7
020FFF9301450F83
00550023FE0F8CE3
5265775300008067
6F53657375462B56
0A736B636F722043
0000000000000000
