0102829300000297
1990006F30529073
00112023FB010113
0041242300312223
0061282300512623
01C12C2300712A23
03E1202301D12E23
02A1242303F12223
02C1282302B12623
02E12C2302D12A23
0501202302F12E23
341022F305112223
300022F304512423
1F0000EF04512623
02051E6300000313
800003B7342022F3
0072F2B3FFF38393
00628A6300B00313
0000009700010513
0410006F13408093
0042829304812283
0900006F04512423
0000339700010293
0043A103D8438393
00512023FF010113
001E0E130003AE03
0003086301C3A023
03C0809300000097
342025730890006F
FFF28293800002B7
158000EF00557533
6EC2829300002297
00A282B300351513
0042A3030002A503
00003317000300E7
00032383D2430313
00732023FFF38393
0002811300012283
02032E0300832383
00003297087E0863
0082A303CFC28293
0293282302832623
03332C2303232A23
0553202303432E23
0573242305632223
0593282305832623
05B32C2305A32A23
0000339702232423
0003AE03B6838393
0202A30307C32623
028321030062A423
0303248302C32403
0383298303432903
04032A8303C32A03
04832B8304432B03
05032C8304C32C03
05832D8305432D03
3412907304812283
3002907304C12283
0041218300012083
00C1228300812203
0141238301012303
01C12E8301812E03
02412F8302012F03
02C1258302812503
0341268303012603
03C1278303812703
0441288304012803
3020007305010113
0000329700000073
0082A303C0C28293
0085751306C32383
00038513300522F3
0010031300008067
3442B37300A312B3
342022F300008067
0062F2B380000337
0002846300000513
0000806700150513
0200079302060063
00F04C6340C787B3
00000713FE060513
0007059300A5D533
00C5D73300008067
00F595B300C55533
FE9FF06F00B56533
0006081300058793
0005031300068893
0000373728069663
0EC5F66384870713
0CD67863000106B7
00C6B6B30FF00693
00D658B300369693
0007470301170733
0200071300D706B3
00070C6340D70733
00D556B300E797B3
00F6E5B300E61833
0108551300E51333
0108161302A5F733
0103569301065613
0107171302A5D5B3
02B607B300D766B3
00F6FE6300058713
FFF58713010686B3
00F6F6630106E863
010686B3FFE58713
02A6F7B340F686B3
0103531301031313
0107979302A6D6B3
02D605B30067E333
00B37C6300068513
FFF6851300680333
00B3746301036663
01071713FFE68513
0000059300A76733
010008B70E40006F
F3166CE301000693
F31FF06F01800693
0010069300061663
000106B702C6D833
0FF006930CD87263
008008930106F463
00D70733011856B3
0200071300074683
40D70733011686B3
410787B30A071863
0108561300100593
0108D89301081893
02C7F73301035693
0107171302C7D7B3
02F8853300D766B3
00A6FE6300078713
FFF78713010686B3
00A6F6630106E863
010686B3FFE78713
02C6F7B340A686B3
0103531301031313
0107979302C6D6B3
02D888B30067E333
01137C6300068513
FFF6851300680333
0113746301036663
01071713FFE68513
0007051300A76733
010006B700008067
F4D862E301000893
F3DFF06F01800893
00D7D5B300E81833
00D556B300E51333
00E797B301085513
00F6E8B302A5F733
0107D79301081793
02A5D5B30108D613
00C7673301071713
0005861302B786B3
0107073300D77E63
01076863FFF58613
FFE5861300D77663
40D706B301070733
0108989302A6F733
02A6D6B30108D893
02D785B301071713
00068713011767B3
010787B300B7FE63
0107E863FFF68713
FFE6871300B7F663
40B787B3010787B3
00E5E5B301061593
18D5E663EB5FF06F
04E6F46300010737
00D837330FF00813
0000383700371713
00E6D5B384880813
0005C803010585B3
00E8083302000593
02059663410585B3
EEF6ECE300100713
0015471300C53533
010005B7EEDFF06F
FCB6E0E301000713
FB9FF06F01800713
00B696B301065733
0106DE9300D766B3
03D778B30107D733
0105583300B797B3
0106979300F86333
010358130107D793
03D7573300B61633
0108E83301089893
00070E1302E78F33
00D8083301E87E63
00D86863FFF70E13
FFE70E1301E87663
41E8083300D80833
03D8583303D878B3
03078EB301089893
0107D79301031793
0008071300F8E7B3
00D787B301D7FE63
00D7E863FFF80713
FFE8071301D7F663
010E1E1300D787B3
00010EB741D787B3
FFFE881300EE6733
0107589301077333
0106561301067833
0308883303030E33
02C30333010E5693
006686B301030333
0106F46302C888B3
0106D61301D888B3
0317E663011608B3
000107B7CF179AE3
00F6F6B3FFF78793
00FE7E3301069693
01C686B300B51533
DAD57CE300000593
CC9FF06FFFF70713
0000071300000593
00003537DA5FF06F
94850513FF010113
0081242300112623
0121202300912223
00452783020010EF
0000061300100693
000005930007A783
0000041300050493
00200913000780E7
0044A783032466B3
0000059300000613
000485130047A783
000780E700140413
0F5010EF3E800513
FF010113FD9FF06F
0081242300112623
02F5046300600793
02050463155010EF
0405166314D010EF
C0058593000035B7
C145051300003537
2D5000EF299000EF
139010EFFFDFF06F
00003437FC051CE3
00842583E3840413
C345051300003537
00842503271000EF
FD1FF06F359010EF
BFC58593000035B7
FB010113FB9FF06F
0491222304812423
0060079304112623
0005841300050493
000037370EA7E063
9507071300251793
0007A78300E787B3
0000353700078067
215000EFA8050513
04442783081010EF
00C4280301042883
0404278302F12823
0004268300442703
03C4278302F12623
0005059304842603
0384278302F12423
B045051300003537
0344278302F12223
0304278302F12023
02C4278300F12E23
0284278300F12C23
0244278300F12A23
0204278300F12823
01C4278300F12623
0184278300F12423
0144278300F12223
0084278300F12023
00040593181000EF
EA9FF0EF00048513
AA85051300003537
00003537F55FF06F
F49FF06FAC450513
0004859300003537
14D000EFAE050513
FF010113F39FF06F
0011262300812423
3420267300050413
0016561300161613
02C7E86300500793
0026179300003737
00F707B396C70713
000035370007A583
105000EF98C50513
0000051300040593
000035B7EA5FF0EF
FE1FF06F98458593
00112623FF010113
00003537342025F3
0015D59300159593
0CD000EFC5C50513
9A858593000035B7
E69FF0EF00400513
D3878793000037B7
00070C630007A703
0007A0230007A303
D3C7A503000037B7
0000806700030067
00112623FF010113
0E5000EF625000EF
0000311767D000EF
000012B7ACC10113
0051013380028293
21C0006FFD9FF0EF
01312E23FD010113
0301268300068993
0321202302812423
0006091300058413
0040061300088593
0211262302912223
00E1262300050493
0101222300F12423
008127830F5010EF
00B405B3FB090593
0604A0230404AE23
02F5A823FF05F593
00C12703000027B7
8807879300412803
000017B704F5A623
0281240302C12083
0335A4239BC78793
0305AA2302E5A623
02B4A42304F5A423
0241248302012903
0301011301C12983
00C0079300008067
00C5278302F58733
00B5070300E787B3
0007A78300B75463
02E6473302000713
0027171301F67513
00F6A02300E787B3
FE01011300008067
00112E2300C10693
00C12703FBDFF0EF
00A7953300100793
01C1208300072783
00F7202300A7E7B3
0000806702010113
0085580300452783
00812423FF010113
0005041302F80833
00A4488300052503
00112623FFF00713
00E405A300912223
00C0031300000593
01F00E1301050533
0315C26302000E93
0084578300000493
00C1208306F4C463
0041248300812403
0000806701010113
00C4260302F85733
00D606B3026586B3
00C6A22300468613
00EE4E6300C6A423
0027D79300B405A3
FFC7F79300378793
FA9FF06F00158593
03D7473301F70713
0027171300A6A023
FD9FF06F00E50533
0004861300442783
02F4873300000593
0004051300042783
00E787B300148493
0047069300C42703
0087268300D7A023
0087268300D7A223
00F7242300F6A023
F51FF06FED5FF0EF
00050793FF010113
0006059300058513
0011262300068613
49C010EF000780E7
00000513718010EF
FF01011300008067
0005041300812423
0011262304500513
0005849300912223
00048593000400E7
000400E705200513
0081240300040313
0004859300C12083
0520051300412483
0003006701010113
001787930005A783
000037B700F5A023
00030067CD07A303
04812423FB010113
03412C2303312E23
0361282303512A23
0491222304112623
0371262305212023
0391222303812423
01B12E2303A12023
00058A9300050A13
00068B1300060993
00E0546300100413
0010079300070413
00FB146302000C13
3B9AD4B703000C13
00A00C9300100913
9FF4849300000713
00A00D1300200D93
0007146300148B93
0379D5330934F263
00190913000A8593
000A00E703050513
FFFC8C9300100713
0379F9B300100793
FCFC96E303A4D4B3
03098513000A8593
00300793000A00E7
06FB0A6341240433
0481240304C12083
0401290304412483
03812A0303C12983
03012B0303412A83
02812C0302C12B83
02012D0302412C83
0501011301C12D83
F9944CE300008067
000A8593F96DEAE3
00E12623000C0513
00190913000A00E7
F79FF06F00C12703
02000513000A8593
FFF40413000A00E7
F8DFF06FFE8048E3
04812423FB010113
0521202304912223
03412C2303312E23
0391222303512A23
01B12E2303A12023
0361282304112623
0381242303712623
0005849300050413
00068D1300060A93
FFF0091300000A13
00000C9300000993
000AC50380000DB7
04C1208304051063
0441248304812403
03C1298304012903
03412A8303812A03
02C12B8303012B03
02412C8302812C03
01C12D8302012D03
0000806705010113
02500693000C9E63
0004859336D50A63
001A8A93000400E7
06400693FA5FF06F
06A6E26310D50E63
02A6EA6303900693
0ED5746303100693
34D50A6302D00693
0CF5006303000793
02E5126302500713
0250051300048593
15C0006F000400E7
1AD50E6305800693
2EE50E6306300713
0250051300048593
00048593000400E7
FD5FF06F000AC503
16D50A6307000693
0690069302A6E063
06C006930AD50263
0680069308D50A63
FC5FF06FF6D506E3
10D5066307500693
0730071302A6EE63
000D2C03FAE518E3
000C0B93004D0B13
26051863000BC503
00F9986300300793
41790BB3418B8BB3
000B0D1327704663
078006930C80006F
07A0069312D50463
00095E63FA9FF06F
FD05091328098863
00200993F00992E3
FE0948E3EFDFF06F
02D9093300A00693
01250933FD090913
001A0A13FE1FF06F
040A1263EDDFF06F
004D0D13000D2603
0004859302065063
00C1202302D00513
00012603000400E7
40C00633FFF90913
0009869300090713
0004051300048593
03C0006FCA1FF0EF
FAEA0EE300100713
FF87F713007D0793
0047268300072603
01B6073300870D13
00D7073300C73733
00048593FA0700E3
C01FF0EF00040513
E59FF06F00000C93
000D2603000A1863
F9DFF06F004D0D13
FEEA08E300100713
FF87F713007D0793
0007260300870D13
FC0710E300472703
FFF7C793800007B7
FB1FF06FF6C7F8E3
0300051300048593
00048593000400E7
000400E707800513
0010099300800913
0B46C26300100693
00012423000D2783
00F12223004D0D13
00000B9301000C13
0100089300012023
0081258300412503
002B1613FFF88B13
9CCFF0EF01112623
0805186300F57513
0300069300012783
00C1288300079863
08F8966300100793
0185151300A68533
4185551300048593
001B8B93000400E7
00300693040B1863
D6D998E300000C93
41770BB300191713
00048593F17054E3
000400E702000513
FEDFF06FFFFB8B93
FF87F693007D0793
00868D130006A783
0046A78300F12223
F55FF06F00F12423
000B089301912023
00900793F59FF06F
F8A7E2E305700693
F7DFF06F03000693
00F12623FFFC0793
0010079301894C63
0004859300F99C63
000400E703000513
FC1FF06F00C12C03
FEF99AE300200793
0200051300048593
00048593FE5FF06F
000400E7001B8B93
00048593D81FF06F
000400E702000513
D85FF06FFFFB8B93
00048593000D2503
000400E7004D0B13
00000A13D75FF06F
00000993FFF00913
C89FF06F00100C93
C81FF06F00300993
C79FF06F00100993
00050613FE010113
0005869300001537
00C10593C5050513
0001262300112E23
01C12083BA1FF0EF
0000806702010113
02B12223FC010113
00112E2302410593
02D1262302C12423
02F12A2302E12823
03112E2303012C23
FA5FF0EF00B12623
0401011301C12083
0000806700008067
3007A7F300800793
0000806710500073
00A7953300100793
0000806730452573
3007B7F300800793
3440507330405073
800017B700008067
0207A5030247A703
FEE59AE30247A583
FE01011300008067
00112E2300812C23
0121282300912A23
0080041301312623
000034B730043473
FC1FF0EFD2848493
0044A9830004A903
4125053300050713
413585B300A73733
090606130003D637
40E585B300000693
0003D7B7FB1FE0EF
02A787B309078793
0127893300847413
013787B300F937B3
00F4A2230124A023
0181240330042473
0141248301C12083
00C1298301012903
2880106F02010113
00112623FF010113
0003D7B7F45FF0EF
8000173709078793
FFF0069300F507B3
00A7B53302D72623
02F7242300B50533
0070051302A72623
00C12083EF1FF0EF
0101011300000513
0C059C6300008067
00812423FF010113
0091222300112623
00050413FFF00793
000047B700F51663
0080049331A78413
ED1FF0EF3004B4F3
FFF4079300004737
0084F49331A70713
0007079308F75463
090705930003D737
000037B702B786B3
0007A603D2878793
08F707930047A803
00A787B340C787B3
3E70071340A60533
02B7D7B300D787B3
00F5053302B787B3
00B787B300A74463
00C7863380001737
02D72623FFF00693
010787B300F637B3
02F7262302C72423
00C120833004A4F3
0041248300812403
0000806701010113
00000793F807D0E3
00008067F79FF06F
00812423FF010113
0080041300112623
E11FF0EF30043473
D287A783000037B7
40F5053300847413
090787930003D7B7
3004247302F55533
0081240300C12083
0000806701010113
0005C70300054783
0007966300E79463
0000806740E78533
0015859300150513
0FF5F693FE1FF06F
0037F71300050793
0FF5F59304071863
00B765B300859713
00B765B301059713
0007871300C78333
40E308B300300813
0026571303186E63
00B787B300271593
02B70733FFC00593
00E7873300C70733
0000806702E79463
00178793FE060EE3
FFF60613FED78FA3
00470713F9DFF06F
FB9FF06FFEB72E23
FED78FA300178793
00852703FD1FF06F
00B7E5B30026F793
04059A6300072503
00C7963300100793
FEA0051300452783
0407806300F677B3
FDD00513F7E6F793
0806F51302079A63
00050A6300472783
00C7222300F66633
0000806700000513
00F67633FFF64613
0000806700C72223
00008067FDD00513
0007A50300852783
000528830047A783
0205906300452803
00C7173300100713
FEA0051300E87833
0006846302080C63
0080071300080693
0008A60330073773
00F647B300877713
0107F7B300D7C7B3
00F8A02300C7C7B3
0000051330072773
0085250300008067
0045250300052703
0007A78300072783
0047250300A7C7B3
0205986300A7F7B3
0017F79300C7D7B3
0010079300F6A023
0047260300C797B3
0007946300C7F7B3
00058513FEA00593
00F6A02300008067
FF1FF06F00000593
0085278300052703
00E7A02300872703
C9078793000037B7
0000051300F52223
0025171300008067
00150513000037B7
00251513CAC78793
00E78733FF010113
0081242300A787B3
0007240300912223
001126230007A483
00C1208300946C63
0041248300812403
0000806701010113
0004051300042783
000780E70047A783
0004222300050463
FCDFF06F00C40413
000037B7FF010113
000034B700912223
0011262300812423
01212023CEC78413
D1048493CEC78793
0005091300941C63
0294146300078413
0440006F00000413
0007086300442703
0007270300042703
00C4041302A70863
00442783FD1FF06F
00C4041300079663
00042783FCDFF06F
0007A58300090513
FE0514E3D21FF0EF
00C1208300040513
0041248300812403
0101011300012903
0000353700008067
D2850613000037B7
40C78633E6478793
D285051300000593
FF010113D05FF06F
0011262300200513
00300513ECDFF0EF
219000EFEC5FF0EF
000037B7EEDFE0EF
00C7C703DC878793
00E78623FFE77713
0101011300C12083
F601011300008067
000047B708812C23
0931262300003437
E3840993C7078793
0101079300F9A223
0000059307000613
08112E2300078513
0921282308912A23
00100713C85FF0EF
0000051300A9A423
E49FF0EF00E10EA3
E41FF0EF00100513
00F11E2310100793
000037B76D0000EF
00003937CC078793
000016B700F12223
000035B700100793
00F12023DC890493
0000079300000713
0000081300000893
400006137DC68693
DC890513E7058593
091000EF0299A023
E384041300D4C783
00E486A3FFB7F713
00079A6301B7F793
000796630184A783
2DC000EFDC890513
CC878793000037B7
0000353700F12223
000026B700100793
D5850493000035B7
00F0089300F12023
0000079300000813
7506869300000713
2705859320000613
021000EFD5850513
0094262300D4C783
FFB7F79300800513
000037B700F486A3
00F42C23E5078793
3005357300F42E23
8BDFE0EF00857513
0005278300452703
00E7A22300F72023
0005222300052023
00D5478300008067
0007986301F7F793
0015351301852503
0000051300008067
FF01011300008067
ABDFF0EF00112623
D4C7A783000037B7
0000373700C12083
E4A7242300A78533
0007851300000593
3990006F01010113
00812423FF010113
0080041300112623
000037B730043473
00950513E407A423
02F5453300A00793
00847413000037B7
000037B7D4A7A623
F91FF0EFD4B7A423
00C1208330042473
0101011300812403
FF01011300008067
0091222300812423
0005049300112623
3004347300800413
00D4C783F21FF0EF
FFD7F79300847413
3004247300F486A3
0081240300C12083
004124830004A423
0000806701010113
E387A783000037B7
0005851300079663
0085F593F98FE06F
000080673005A5F3
E387270300003737
F7CFE06F00071463
3007A7F300857793
0080051300008067
0085751330053573
00800793FD9FF06F
000037373007B7F3
00F6C703E4072683
00E687A3FFF70713
3007A7F30087F793
0005278300008067
0000079300F51463
0000806700078513
00812C23FE010113
00912A2300003437
E384051300050493
00112E2302450513
E3840413FCDFF0EF
00C4250300051463
02049A6300842783
01F7771300D7C703
00E7D68302071463
00D77E6307F00713
01C1208302F42023
0141248301812403
0000806702010113
00A1262300F50863
00C12503E35FF0EF
FD9FF06F02A42023
00812423FF010113
0080041300112623
000037B730043473
00100513E407A703
00F7478300847413
00F707A300178793
30042473F51FF0EF
00C1208300812403
EF1FF06F01010113
00812423FF010113
0080041300112623
0000373730043473
0247A783E3870793
E5C68693000036B7
E387071300847413
04078E6306D78063
00E5060302872583
0506506300E78803
00F520230047A703
00A7202300E52223
00D5478300A7A223
00F506A30407E793
ECDFF0EF00000513
00C1208330042473
0101011300812403
00B7866300008067
FA079AE30007A783
00D5202302872783
0287278300F52223
02A7242300A7A023
FF052783FB5FF06F
00812423FF010113
0011262301212023
0005041300912223
02078663FE850913
3004B4F300800493
CC5FF0EF00090513
0084F493FF544783
FEF40AA3FFD7F793
FE0428233004A4F3
00090513FF544783
FEF40AA3FEB7F793
02050063CB5FF0EF
00C1208300812403
0009051300412483
0101011300012903
00C12083ED9FF06F
0041248300812403
0101011300012903
FF01011300008067
0091222300812423
0005041300112623
3004B4F300800493
00003737C41FF0EF
0247A783E3870793
E5C68693000036B7
E38707130084F493
0607846306D78663
00E4060302872583
04A6566300E78503
00F420230047A683
0086A02300D42223
00D447830087A223
0407E79300872503
00F406A340850533
D75FF0EF00153513
00C120833004A4F3
0041248300812403
0000806701010113
0007A78300B78663
02872783FA0794E3
00F4222300D42023
0087A02302872783
FA9FF06F02872423
D4C7A783000037B7
000037B706078663
0087A703E3878793
00E7560307F00693
000036B704C6EA63
D486A68300E70603
000036B704D64263
02D70C63CE86A683
0206986301872683
02D540630107A683
00070513FF010113
EE1FF0EF00112623
0101011300C12083
40A686B3B6DFF06F
0000806700D7A823
00812423FF010113
0011262300912223
0080041300050493
00D5478330043473
0407F79300847413
AF5FF0EF00078A63
FBF7F79300D4C783
000037B700F486A3
40950533E407A503
C6DFF0EF00153513
00C1208330042473
0041248300812403
0000806701010113
00812C23FE010113
0131262301212823
0015099300112E23
065000EF00912A23
0080091300A98433
000034B730093973
0084A503E3848493
0084A503F61FF0EF
00098613000025B7
01850513C7C58593
0084A703518000EF
00D7478300897513
00F706A30107E793
015000EFB08FE0EF
0005546340A40533
01C1208300000513
0141248301812403
00C1298301012903
0000806702010113
E3878793000037B7
02E7A22302478713
0000059302E7A423
A75FF06F00000513
00812423FF010113
E384079300003437
000037B70087A703
00112623CE87A783
06F7026300912223
00800493E3840413
008425033004B4F3
9C5FF0EF0084F493
000036B702442783
00842703E5C68693
0607806306D78263
00E7058302842603
04A5D26300E78503
00F720230047A683
00E6A02300D72223
0010051300E7A223
3004A4F3B19FF0EF
3005357300800513
00C1208300812403
0085751300412483
A14FE06F01010113
0007A78300F60663
02842783FA0798E3
00F7222300D72023
00E7A02302842783
FB1FF06F02E42423
00A0079300950513
FE01011302F54533
02051A6300112E23
F15FF0EF00A12623
3E80079300C12503
0640061302F515B3
02F5053300000693
01C12083A38FE0EF
0000806702010113
FD9FF06FE31FF0EF
E407A503000037B7
00D5478300008067
0007986301F7F793
0015351301852503
0000051300008067
000037B700008067
00A03533E387A503
000037B700008067
00C7C503E407A783
0000806700157513
00812423FF010113
0091222300112623
3004347300800413
0084741300D54783
00071E630047F713
00C1208330042473
0041248300812403
0000806701010113
00F506A3FFB7F793
F71FF0EF00050493
0004851300050663
00040593A99FF0EF
00C1208300812403
0000353700412483
01010113E6450513
FE010113929FF06F
00812C2302012303
0061202300112E23
84DFE0EF00050413
E407A783000037B7
0687A78301C12083
0181240306F42423
0000806702010113
FF01011306052783
0011262300812423
0007846300050413
00040513000780E7
02050463EE5FF0EF
C8DFF0EF00040513
00C1208300D44783
00F406A30087E793
0101011300812403
00D4478300008067
000786630027F793
841FF0EF00040513
FC0786E301842783
2FC000EF01840513
FD010113FC1FF06F
03212023000037B7
0281242300003937
0211262302912223
01412C2301312E23
D1078493D1078413
03246E63D1090913
889FF0EF00048413
00A00993FFF00493
0724646300002A37
02C1208302812403
0201290302412483
01812A0301C12983
915FF06F03010113
00F1222302C42783
00F1202302042783
01C4288301442783
0104270301842803
0084260300C42683
0004250300442583
00042783EB5FF0EF
030404130487AE23
02442603F85FF06F
0004250300960863
E15FF0EF00061863
F81FF06F03040413
0336463300960613
01850513C7CA0593
134000EF00160613
00D50623FE1FF06F
00B5072300C506A3
00052C23000507A3
0000806700052E23
02112623FD010113
3005B5F300800593
00B126230085F593
00C12583E71FF0EF
F4CFF0EF01C10513
0301011302C12083
000037B700008067
00079463D507A783
00000513920FF06F
0005278300008067
0000373702050263
00E50C63CD872703
0087A70300078A63
00D7073300852683
0045270300E7A423
00E7A22300F72023
0005222300052023
000037B700008067
FF010113D547C783
0081242300112623
FFF0051300912223
8000053700079663
000037B7FFF54513
0007A403CD478793
0204026302F40463
F69FF0EF00842483
0000051340A484B3
008424030004C863
40A40533F55FF0EF
E487A783000037B7
00A7D46300078663
00C1208300078513
0041248300812403
0000806701010113
00812C23FE010113
00112E2300912A23
00C1262300050413
0080049300B52623
F01FF0EF3004B4F3
0084F49300C12603
0010061300C04463
CD47A703000037B7
00C4242300A60633
00F70663CD478793
020710630047A583
00F420230047A703
0047A70300E42223
0087A22300872023
0087260302C0006F
04C6D86300842683
00D7242340D606B3
00E4202300472683
0086A02300D42223
0007A70300872223
00E4186300F70A63
00000593ED5FF0EF
3004A4F3EC5FE0EF
0181240301C12083
0201011301412483
40C686B300008067
F8B702E300D42423
F79FF06F00072703
00812423FF010113
0080041300112623
0005278330043473
0207806300847413
00000513E3DFF0EF
00C1208330042473
0101011300812403
FEA0051300008067
FF010113FE9FF06F
0081242300112623
3007B47300800793
00847793E45FF0EF
00C120833007A7F3
0101011300812403
FE01011300008067
00912A2300812C23
0005049300112E23
0080041300B12623
E09FF0EF30043473
00C1258300847413
0010079300A4DA63
0004851300A7D663
30042473DE5FE0EF
0181240301C12083
0201011301412483
FE01011300008067
00912A2300812C23
0121282300112E23
0141242301312623
0005049301512223
FE4FF0EF00800413
000039B730043473
0000393700003A37
00847413D499A823
CD4A0A13D5098993
00800A93D3090913
0009A783000A2483
0049250300092683
00048A6301448C63
06E7D0630084A703
00E4A42340F70733
41F7D71300D786B3
00F6B7B300A70733
00D9202300E787B3
0009A02300F92223
00000593D35FF0EF
30042473D25FE0EF
0181240301C12083
0101290301412483
00812A0300C12983
0201011300412A83
00D706B300008067
00A585B341F75593
00B6063300E6B633
0004A42340E787B3
00D9202300048513
00F9A02300C92223
30042473C95FF0EF
0004851300C4A783
300AB473000780E7
F3DFF06F00847413
00812423FF010113
0080041300112623
D75FE0EF30043473
D307071300003737
0007250300050793
0084741300472583
00F537B300A78533
3004247300B785B3
0081240300C12083
0000806701010113
00112623FF010113
00C12083FA9FF0EF
0000806701010113
00812423FF010113
0011262300912223
0020049300800413
DD9FF0EF300437F3
0010051300A4C463
DF9FF0EF00100593
FE5FF06FAE1FE0EF
00812423FF010113
0000343700912223
00112623000034B7
D1048493D1040413
00C1208300946E63
0041248300812403
0101011300000513
0144079300008067
00F42A2300040513
B04FE0EF00F42C23
FCDFF06F01C40413
0000000000008067
0000000000000938
0000000000000938
0000000000000938
0000000000000938
0000000000000938
0000000000000938
0000000000000938
00002948000012AC
00002CDC00001690
0000134800002C84
000029A400000000
0000000000002788
0303030302020100
0404040404040404
0505050505050505
0505050505050505
0606060606060606
0606060606060606
0606060606060606
0606060606060606
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
000000003044454C
000008C800000810
00000804000008C8
000008B000000810
000029F8000008BC
00002A3400002A18
00002A5400002A48
6E6B6E7500002A6C
65637845006E776F
6163206E6F697470
2820732520657375
000000000A296425
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
7463757274736E49
72646461206E6F69
6173696D20737365
000064656E67696C
7463757274736E49
65636341206E6F69
746C756166207373
656C6C4900000000
74736E69206C6167
006E6F6974637572
696F706B61657242
64616F4C0000746E
7373657264646120
67696C6173696D20
64616F4C0064656E
2073736563636120
000000746C756166
72654B202A2A2A2A
6F6C6C41206C656E
46206E6F69746163
20216572756C6961
0000000A2A2A2A2A
654B202A2A2A2A2A
504F4F206C656E72
2A2A2A2A2A202153
2A2A2A2A0000000A
6C656E72654B202A
202163696E615020
00000A2A2A2A2A2A
6B6E55202A2A2A2A
746146206E776F6E
726F727245206C61
2A2A2A2021642520
7272754300000A2A
6572687420746E65
203D204449206461
746C7561460A7025
74736E6920676E69
206E6F6974637572
2073736572646461
200A78257830203D
257830203A617220
30203A7067202078
3A70742020782578
7420207825783020
0A78257830203A30
7830203A31742020
203A327420207825
3374202078257830
202078257830203A
78257830203A3474
30203A357420200A
3A36742020782578
6120207825783020
2078257830203A30
257830203A316120
203A326120200A78
3361202078257830
202078257830203A
78257830203A3461
7830203A35612020
3A366120200A7825
6120207825783020
0A78257830203A37
0052534900000000
6169746E65737365
646165726874206C
6174614600000000
20746C756166206C
5320217325206E69
2E676E696E6E6970
61746146000A2E2E
20746C756166206C
6165726874206E69
6241202170252064
0A2E676E6974726F
7275705300000000
746E692073756F69
6420747075727265
2164657463657465
6425203A51524920
5F7379730000000A
0000006B636F6C63
000015D000001564
0000000000001634
0000000000000000
00002CEC00000000
00002D1000002D04
00002D1000002D10
000000006E69616D
FFFFFF00656C6469
00002CD400000BFC
8000101000002CD4
FFFFFFF500000001
0000283C00002D58
0000000000000000
0000000000002824
0000283000002D40
0000000000000000
00002D1000002D10
0000000000000000
000000000000000F
