000073B32BC00313
FE731EE300138393
00A3031380001337
FE038EE300034383
04018193800011B7
0201802300300993
041003130FF0000F
0FF0000F00618023
0261802300100313
003005130FF0000F
0C0000EF0C4000EF
08098263FFF98993
5273031356190337
0A8000EFFCB312E3
0A0000EF0A4000EF
0006041306C000EF
060000EF094000EF
088000EF00060493
00060913054000EF
078000EF07C000EF
070000EF074000EF
068000EF06C000EF
060000EF064000EF
058000EF05C000EF
050000EF00000A13
00B3202301448333
004A0A130FF0000F
00090067FF4456E3
018596130000006F
0FF373130085D313
0066663301031313
0FF373130105D313
0066663300831313
006666330185D313
0040029300008067
0FF0000F00A18823
0FF0000F0081C303
FE031AE300137313
0101C3030085D593
0065E5B301831313
FFF2829300855513
00008067FC0298E3
0000000000000000
