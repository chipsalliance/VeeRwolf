7C029073AAAA02B7
00000797098000EF
0D0000EF0FC78793
00A3031380001337
FE038EE300034383
0F67879300000797
800013370B4000EF
0023538301030313
00000E1300E3D393
001E0E1303C38263
001E0E1303C38663
0000079703C38A63
080000EF10D78793
000007970340006F
070000EF0BB78793
000007971080006F
060000EF0C478793
000007972380006F
050000EF0CA78793
0000006F00000067
08000E1380002737
80001E3701C70623
000E2E8303CE0E13
200E0E130001CE37
004E5E9303CEDE33
00300E1301D70023
08700E1301C70623
0007022301C70423
0007828300008067
020FFF9301470F83
00570023FE0F8CE3
0007828300178793
00008067FE0294E3
20676E69746F6F42
666C6F5652657753
4152000A0D2E2E2E
42000A0D4B4F204D
6620676E69746F6F
20495053206D6F72
000A0D6873616C46
20676E69746F6F42
726573206D6F7266
6F42000A0D6C6169
726620676E69746F
0A0D4D4152206D6F
6E776F6E6B6E5500
6F6D20746F6F6220
000000000A0D6564
000073B32BC00313
FE731EE300138393
04018193800011B7
0201802300300993
041003130FF0000F
0FF0000F00618023
0261802300100313
003005130FF0000F
0C0000EF0C4000EF
00099463FFF98993
56190337ECDFF06F
FCB310E352730313
0A0000EF0A4000EF
068000EF09C000EF
090000EF00060413
0006049305C000EF
050000EF084000EF
078000EF00060913
070000EF074000EF
068000EF06C000EF
060000EF064000EF
058000EF05C000EF
00000A13054000EF
0144833304C000EF
0FF0000F00B32023
FF4456E3004A0A13
0185961300090067
0FF373130085D313
0066663301031313
0FF373130105D313
0066663300831313
006666330185D313
0040029300008067
0FF0000F00A18823
0FF0000F0081C303
FE031AE300137313
0101C3030085D593
0065E5B301831313
FFF2829300855513
00008067FC0298E3
00000F9300000F13
0000019300000613
00058E03800025B7
0000043303A00313
FE651EE30F0002EF
088000EF001F8F93
080000EF00050213
078000EF00851113
070000EF00A16133
FFF5051302050C63
0940006F00050463
01E5802304700F13
06F00F130FF0000F
0FF0000F01E58023
01E5802302100F13
000600670FF0000F
0041023300218133
00A1002302C000EF
FE221AE300110113
0FF4741301C000EF
02E00F1304041463
0FF0000F01E58023
05C002EFF71FF06F
FF95051300654463
00451393FD050513
00654463048002EF
FD050513FF950513
0FF5751300756533
0000806700A40433
01E5802304500F13
01E5802307200F13
06F00F1301E58023
07200F1301E58023
FDDFF06F01E58023
0015751301458503
00058503FE050CE3
0000000000028067
