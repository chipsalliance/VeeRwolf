0105051380001537
0010031300255283
000384630012F393
0012D29300131313
FFF30313FE0298E3
FD5FF06F00651023
0000000000000000
