// SPDX-License-Identifier: Apache-2.0
// Copyright 2019 Western Digital Corporation or its affiliates.
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

//********************************************************************************
// $Id$
//
// Function: SweRVolf tech-agnostic toplevel
// Comments:
//
//********************************************************************************

`default_nettype none
module swervolf_core
  #(parameter bootrom_file  = "")
   (input wire 	clk,
    input wire 	       rstn,
    input wire 	       dmi_reg_en,
    input wire [6:0]   dmi_reg_addr,
    input wire 	       dmi_reg_wr_en,
    input wire [31:0]  dmi_reg_wdata,
    output wire [31:0] dmi_reg_rdata,
    input wire 	       dmi_hard_reset,
    output wire        o_flash_sclk,
    output wire        o_flash_cs_n,
    output wire        o_flash_mosi,
    input wire 	       i_flash_miso,
    output wire        o_sd_sclk,
    output wire        o_sd_cs_n,
    output wire        o_sd_mosi,
    input wire 	       i_sd_miso,
    input wire 	       i_uart_rx,
    output wire        o_uart_tx,
    input wire         i_ethmac_mtx_clk,
    output wire [3:0]  o_ethmac_mtxd,
    output wire        o_ethmac_mtxen,
    output wire        o_ethmac_mtxerr,
    input wire         i_ethmac_mrx_clk,
    input wire  [3:0]  i_ethmac_mrxd,
    input wire         i_ethmac_mrxdv,
    input wire         i_ethmac_mrxerr,
    input wire         i_ethmac_mcoll,
    input wire         i_ethmac_mcrs,
    output wire        o_ethmac_mdc,
    input wire         i_ethmac_md,
    output wire        o_ethmac_md,
    output wire        o_ethmac_mdoe,
    output wire [5:0]  o_ram_awid,
    output wire [31:0] o_ram_awaddr,
    output wire [7:0]  o_ram_awlen,
    output wire [2:0]  o_ram_awsize,
    output wire [1:0]  o_ram_awburst,
    output wire        o_ram_awlock,
    output wire [3:0]  o_ram_awcache,
    output wire [2:0]  o_ram_awprot,
    output wire [3:0]  o_ram_awregion,
    output wire [3:0]  o_ram_awqos,
    output wire        o_ram_awvalid,
    input wire 	       i_ram_awready,
    output wire [5:0]  o_ram_arid,
    output wire [31:0] o_ram_araddr,
    output wire [7:0]  o_ram_arlen,
    output wire [2:0]  o_ram_arsize,
    output wire [1:0]  o_ram_arburst,
    output wire        o_ram_arlock,
    output wire [3:0]  o_ram_arcache,
    output wire [2:0]  o_ram_arprot,
    output wire [3:0]  o_ram_arregion,
    output wire [3:0]  o_ram_arqos,
    output wire        o_ram_arvalid,
    input wire 	       i_ram_arready,
    output wire [63:0] o_ram_wdata,
    output wire [7:0]  o_ram_wstrb,
    output wire        o_ram_wlast,
    output wire        o_ram_wvalid,
    input wire 	       i_ram_wready,
    input wire [5:0]   i_ram_bid,
    input wire [1:0]   i_ram_bresp,
    input wire 	       i_ram_bvalid,
    output wire        o_ram_bready,
    input wire [5:0]   i_ram_rid,
    input wire [63:0]  i_ram_rdata,
    input wire [1:0]   i_ram_rresp,
    input wire 	       i_ram_rlast,
    input wire 	       i_ram_rvalid,
    output wire        o_ram_rready,
    input wire 	       i_ram_init_done,
    input wire 	       i_ram_init_error,
    output wire        o_gpio);

   localparam BOOTROM_SIZE = 32'h1000;

   wire        rst_n = rstn;
   wire        timer_irq;
   wire        uart_irq;
   wire        spi0_irq;
   wire        spi1_irq;
   wire        ethmac_irq;

`include "axi_intercon.vh"

   assign o_ram_awid     = ram_awid;
   assign o_ram_awaddr   = ram_awaddr;
   assign o_ram_awlen    = ram_awlen;
   assign o_ram_awsize   = ram_awsize;
   assign o_ram_awburst  = ram_awburst;
   assign o_ram_awlock   = ram_awlock;
   assign o_ram_awcache  = ram_awcache;
   assign o_ram_awprot   = ram_awprot;
   assign o_ram_awregion = ram_awregion;
   assign o_ram_awqos    = ram_awqos;
   assign o_ram_awvalid  = ram_awvalid;
   assign ram_awready    = i_ram_awready;
   assign o_ram_arid     = ram_arid;
   assign o_ram_araddr   = ram_araddr;
   assign o_ram_arlen    = ram_arlen;
   assign o_ram_arsize   = ram_arsize;
   assign o_ram_arburst  = ram_arburst;
   assign o_ram_arlock   = ram_arlock;
   assign o_ram_arcache  = ram_arcache;
   assign o_ram_arprot   = ram_arprot;
   assign o_ram_arregion = ram_arregion;
   assign o_ram_arqos    = ram_arqos;
   assign o_ram_arvalid  = ram_arvalid;
   assign ram_arready    = i_ram_arready;
   assign o_ram_wdata    = ram_wdata;
   assign o_ram_wstrb    = ram_wstrb;
   assign o_ram_wlast    = ram_wlast;
   assign o_ram_wvalid   = ram_wvalid;
   assign ram_wready     = i_ram_wready;
   assign ram_bid        = i_ram_bid;
   assign ram_bresp      = i_ram_bresp;
   assign ram_bvalid     = i_ram_bvalid;
   assign o_ram_bready   = ram_bready;
   assign ram_rid        = i_ram_rid;
   assign ram_rdata      = i_ram_rdata;
   assign ram_rresp      = i_ram_rresp;
   assign ram_rlast      = i_ram_rlast;
   assign ram_rvalid     = i_ram_rvalid;
   assign o_ram_rready   = ram_rready;

   axi_mem_wrapper
     #(.ID_WIDTH  (`RV_LSU_BUS_TAG+2),
       .MEM_SIZE  (BOOTROM_SIZE),
       .INIT_FILE (bootrom_file))
   bootrom
     (.clk      (clk),
      .rst_n    (rst_n),
      .i_awid    (rom_awid),
      .i_awaddr  (rom_awaddr),
      .i_awlen   (rom_awlen),
      .i_awsize  (rom_awsize),
      .i_awburst (rom_awburst),
      .i_awvalid (rom_awvalid),
      .o_awready (rom_awready),

      .i_arid    (rom_arid),
      .i_araddr  (rom_araddr),
      .i_arlen   (rom_arlen),
      .i_arsize  (rom_arsize),
      .i_arburst (rom_arburst),
      .i_arvalid (rom_arvalid),
      .o_arready (rom_arready),

      .i_wdata  (rom_wdata),
      .i_wstrb  (rom_wstrb),
      .i_wlast  (rom_wlast),
      .i_wvalid (rom_wvalid),
      .o_wready (rom_wready),

      .o_bid    (rom_bid),
      .o_bresp  (rom_bresp),
      .o_bvalid (rom_bvalid),
      .i_bready (rom_bready),

      .o_rid    (rom_rid),
      .o_rdata  (rom_rdata),
      .o_rresp  (rom_rresp),
      .o_rlast  (rom_rlast),
      .o_rvalid (rom_rvalid),
      .i_rready (rom_rready));

   axi_multicon
     #(.ID_WIDTH  (`RV_LSU_BUS_TAG+2))
   multicon
     (.clk       (clk),
      .rst_n     (rst_n),
      .o_gpio    (o_gpio),
      .o_sclk0   (o_flash_sclk),
      .o_cs_n0   (o_flash_cs_n),
      .o_mosi0   (o_flash_mosi),
      .i_miso0   (i_flash_miso),
      .o_sclk1   (o_sd_sclk),
      .o_cs_n1   (o_sd_cs_n),
      .o_mosi1   (o_sd_mosi),
      .i_miso1   (i_sd_miso),
      .o_spi0_irq  (spi0_irq),
      .o_spi1_irq  (spi1_irq),
      .o_timer_irq (timer_irq),
      .i_ram_init_done  (i_ram_init_done),
      .i_ram_init_error (i_ram_init_error),
      .i_awid    (multicon_awid),
      .i_awaddr  (multicon_awaddr),
      .i_awlen   (multicon_awlen),
      .i_awsize  (multicon_awsize),
      .i_awburst (multicon_awburst),
      .i_awvalid (multicon_awvalid),
      .o_awready (multicon_awready),
      .i_arid    (multicon_arid),
      .i_araddr  (multicon_araddr),
      .i_arlen   (multicon_arlen),
      .i_arsize  (multicon_arsize),
      .i_arburst (multicon_arburst),
      .i_arvalid (multicon_arvalid),
      .o_arready (multicon_arready),
      .i_wdata   (multicon_wdata),
      .i_wstrb   (multicon_wstrb),
      .i_wlast   (multicon_wlast),
      .i_wvalid  (multicon_wvalid),
      .o_wready  (multicon_wready),
      .o_bid     (multicon_bid),
      .o_bresp   (multicon_bresp),
      .o_bvalid  (multicon_bvalid),
      .i_bready  (multicon_bready),
      .o_rid     (multicon_rid),
      .o_rdata   (multicon_rdata),
      .o_rresp   (multicon_rresp),
      .o_rlast   (multicon_rlast),
      .o_rvalid  (multicon_rvalid),
      .i_rready  (multicon_rready));

   axi_uart_wrapper
     #(.ID_WIDTH  (`RV_LSU_BUS_TAG+2))
   uart
     (.clk        (clk),
      .rst_n      (rst_n),
      .i_uart_rx  (i_uart_rx),
      .o_uart_tx  (o_uart_tx),
      .o_uart_irq (uart_irq),
      .i_awid     (uart_awid),
      .i_awaddr   (uart_awaddr[11:0]),
      .i_awlen    (uart_awlen),
      .i_awsize   (uart_awsize),
      .i_awburst  (uart_awburst),
      .i_awvalid  (uart_awvalid),
      .o_awready  (uart_awready),
      .i_arid     (uart_arid),
      .i_araddr   (uart_araddr[11:0]),
      .i_arlen    (uart_arlen),
      .i_arsize   (uart_arsize),
      .i_arburst  (uart_arburst),
      .i_arvalid  (uart_arvalid),
      .o_arready  (uart_arready),
      .i_wdata    (uart_wdata),
      .i_wstrb    (uart_wstrb),
      .i_wlast    (uart_wlast),
      .i_wvalid   (uart_wvalid),
      .o_wready   (uart_wready),
      .o_bid      (uart_bid),
      .o_bresp    (uart_bresp),
      .o_bvalid   (uart_bvalid),
      .i_bready   (uart_bready),
      .o_rid      (uart_rid),
      .o_rdata    (uart_rdata),
      .o_rresp    (uart_rresp),
      .o_rlast    (uart_rlast),
      .o_rvalid   (uart_rvalid),
      .i_rready   (uart_rready));

   axi_ethmac_wrapper
     #(.ID_WIDTH  (`RV_LSU_BUS_TAG+2))
   ethmac
     (.clk          (clk),
      .rst_n        (rst_n),
      .o_dma_awid     (ethmac_dma_awid    ),
      .o_dma_awaddr   (ethmac_dma_awaddr  ),
      .o_dma_awlen    (ethmac_dma_awlen   ),
      .o_dma_awsize   (ethmac_dma_awsize  ),
      .o_dma_awburst  (ethmac_dma_awburst ),
      .o_dma_awlock   (ethmac_dma_awlock  ),
      .o_dma_awcache  (ethmac_dma_awcache ),
      .o_dma_awprot   (ethmac_dma_awprot  ),
      .o_dma_awregion (ethmac_dma_awregion),
      .o_dma_awqos    (ethmac_dma_awqos   ),
      .o_dma_awvalid  (ethmac_dma_awvalid ),
      .i_dma_awready  (ethmac_dma_awready ),
      .o_dma_arid     (ethmac_dma_arid    ),
      .o_dma_araddr   (ethmac_dma_araddr  ),
      .o_dma_arlen    (ethmac_dma_arlen   ),
      .o_dma_arsize   (ethmac_dma_arsize  ),
      .o_dma_arburst  (ethmac_dma_arburst ),
      .o_dma_arlock   (ethmac_dma_arlock  ),
      .o_dma_arcache  (ethmac_dma_arcache ),
      .o_dma_arprot   (ethmac_dma_arprot  ),
      .o_dma_arregion (ethmac_dma_arregion),
      .o_dma_arqos    (ethmac_dma_arqos   ),
      .o_dma_arvalid  (ethmac_dma_arvalid ),
      .i_dma_arready  (ethmac_dma_arready ),
      .o_dma_wdata    (ethmac_dma_wdata   ),
      .o_dma_wstrb    (ethmac_dma_wstrb   ),
      .o_dma_wlast    (ethmac_dma_wlast   ),
      .o_dma_wvalid   (ethmac_dma_wvalid  ),
      .i_dma_wready   (ethmac_dma_wready  ),
      .i_dma_bid      (ethmac_dma_bid     ),
      .i_dma_bresp    (ethmac_dma_bresp   ),
      .i_dma_bvalid   (ethmac_dma_bvalid  ),
      .o_dma_bready   (ethmac_dma_bready  ),
      .i_dma_rid      (ethmac_dma_rid     ),
      .i_dma_rdata    (ethmac_dma_rdata   ),
      .i_dma_rresp    (ethmac_dma_rresp   ),
      .i_dma_rlast    (ethmac_dma_rlast   ),
      .i_dma_rvalid   (ethmac_dma_rvalid  ),
      .o_dma_rready   (ethmac_dma_rready  ),
      .i_awid     (ethmac_awid),
      .i_awaddr   (ethmac_awaddr[11:0]),
      .i_awlen    (ethmac_awlen),
      .i_awsize   (ethmac_awsize),
      .i_awburst  (ethmac_awburst),
      .i_awvalid  (ethmac_awvalid),
      .o_awready  (ethmac_awready),
      .i_arid     (ethmac_arid),
      .i_araddr   (ethmac_araddr[11:0]),
      .i_arlen    (ethmac_arlen),
      .i_arsize   (ethmac_arsize),
      .i_arburst  (ethmac_arburst),
      .i_arvalid  (ethmac_arvalid),
      .o_arready  (ethmac_arready),
      .i_wdata    (ethmac_wdata),
      .i_wstrb    (ethmac_wstrb),
      .i_wlast    (ethmac_wlast),
      .i_wvalid   (ethmac_wvalid),
      .o_wready   (ethmac_wready),
      .o_bid      (ethmac_bid),
      .o_bresp    (ethmac_bresp),
      .o_bvalid   (ethmac_bvalid),
      .i_bready   (ethmac_bready),
      .o_rid      (ethmac_rid),
      .o_rdata    (ethmac_rdata),
      .o_rresp    (ethmac_rresp),
      .o_rlast    (ethmac_rlast),
      .o_rvalid   (ethmac_rvalid),
      .i_rready   (ethmac_rready),
      .i_mtx_clk_pad (i_ethmac_mtx_clk),
      .o_mtxd_pad    (o_ethmac_mtxd),
      .o_mtxen_pad   (o_ethmac_mtxen),
      .o_mtxerr_pad  (o_ethmac_mtxerr),
      .i_mrx_clk_pad (i_ethmac_mrx_clk),
      .i_mrxd_pad    (i_ethmac_mrxd),
      .i_mrxdv_pad   (i_ethmac_mrxdv),
      .i_mrxerr_pad  (i_ethmac_mrxerr),
      .i_mcoll_pad   (i_ethmac_mcoll),
      .i_mcrs_pad    (i_ethmac_mcrs),
      .o_mdc_pad     (o_ethmac_mdc),
      .i_md_pad      (i_ethmac_md),
      .o_md_pad      (o_ethmac_md),
      .o_md_padoe    (o_ethmac_mdoe),
      .o_int         (ethmac_irq)
      );


   swerv_wrapper_dmi rvtop
     (
      .clk     (clk),
      .rst_l   (rstn),
      .rst_vec (31'h40000000),
      .nmi_int (1'b0),
      .nmi_vec (31'h8880000),

      .trace_rv_i_insn_ip      (),
      .trace_rv_i_address_ip   (),
      .trace_rv_i_valid_ip     (),
      .trace_rv_i_exception_ip (),
      .trace_rv_i_ecause_ip    (),
      .trace_rv_i_interrupt_ip (),
      .trace_rv_i_tval_ip      (),

      // Bus signals
      //-------------------------- LSU AXI signals--------------------------
      .lsu_axi_awvalid  (lsu_awvalid),
      .lsu_axi_awready  (lsu_awready),
      .lsu_axi_awid     (lsu_awid   ),
      .lsu_axi_awaddr   (lsu_awaddr ),
      .lsu_axi_awregion (lsu_awregion),
      .lsu_axi_awlen    (lsu_awlen  ),
      .lsu_axi_awsize   (lsu_awsize ),
      .lsu_axi_awburst  (lsu_awburst),
      .lsu_axi_awlock   (lsu_awlock ),
      .lsu_axi_awcache  (lsu_awcache),
      .lsu_axi_awprot   (lsu_awprot ),
      .lsu_axi_awqos    (lsu_awqos  ),

      .lsu_axi_wvalid   (lsu_wvalid),
      .lsu_axi_wready   (lsu_wready),
      .lsu_axi_wdata    (lsu_wdata),
      .lsu_axi_wstrb    (lsu_wstrb),
      .lsu_axi_wlast    (lsu_wlast),

      .lsu_axi_bvalid   (lsu_bvalid),
      .lsu_axi_bready   (lsu_bready),
      .lsu_axi_bresp    (lsu_bresp ),
      .lsu_axi_bid      (lsu_bid   ),

      .lsu_axi_arvalid  (lsu_arvalid ),
      .lsu_axi_arready  (lsu_arready ),
      .lsu_axi_arid     (lsu_arid    ),
      .lsu_axi_araddr   (lsu_araddr  ),
      .lsu_axi_arregion (lsu_arregion),
      .lsu_axi_arlen    (lsu_arlen   ),
      .lsu_axi_arsize   (lsu_arsize  ),
      .lsu_axi_arburst  (lsu_arburst ),
      .lsu_axi_arlock   (lsu_arlock  ),
      .lsu_axi_arcache  (lsu_arcache ),
      .lsu_axi_arprot   (lsu_arprot  ),
      .lsu_axi_arqos    (lsu_arqos   ),

      .lsu_axi_rvalid   (lsu_rvalid),
      .lsu_axi_rready   (lsu_rready),
      .lsu_axi_rid      (lsu_rid   ),
      .lsu_axi_rdata    (lsu_rdata ),
      .lsu_axi_rresp    (lsu_rresp ),
      .lsu_axi_rlast    (lsu_rlast ),

      //-------------------------- IFU AXI signals--------------------------
      .ifu_axi_awvalid  (),
      .ifu_axi_awready  (1'b0),
      .ifu_axi_awid     (),
      .ifu_axi_awaddr   (),
      .ifu_axi_awregion (),
      .ifu_axi_awlen    (),
      .ifu_axi_awsize   (),
      .ifu_axi_awburst  (),
      .ifu_axi_awlock   (),
      .ifu_axi_awcache  (),
      .ifu_axi_awprot   (),
      .ifu_axi_awqos    (),

      .ifu_axi_wvalid   (),
      .ifu_axi_wready   (1'b0),
      .ifu_axi_wdata    (),
      .ifu_axi_wstrb    (),
      .ifu_axi_wlast    (),

      .ifu_axi_bvalid   (1'b0),
      .ifu_axi_bready   (),
      .ifu_axi_bresp    (2'b00),
      .ifu_axi_bid      (3'd0),

      .ifu_axi_arvalid  (ifu_arvalid ),
      .ifu_axi_arready  (ifu_arready ),
      .ifu_axi_arid     (ifu_arid    ),
      .ifu_axi_araddr   (ifu_araddr  ),
      .ifu_axi_arregion (ifu_arregion),
      .ifu_axi_arlen    (ifu_arlen   ),
      .ifu_axi_arsize   (ifu_arsize  ),
      .ifu_axi_arburst  (ifu_arburst ),
      .ifu_axi_arlock   (ifu_arlock  ),
      .ifu_axi_arcache  (ifu_arcache ),
      .ifu_axi_arprot   (ifu_arprot  ),
      .ifu_axi_arqos    (ifu_arqos   ),

      .ifu_axi_rvalid   (ifu_rvalid),
      .ifu_axi_rready   (ifu_rready),
      .ifu_axi_rid      (ifu_rid   ),
      .ifu_axi_rdata    (ifu_rdata ),
      .ifu_axi_rresp    (ifu_rresp ),
      .ifu_axi_rlast    (ifu_rlast ),

      //-------------------------- SB AXI signals-------------------------
      .sb_axi_awvalid  (sb_awvalid ),
      .sb_axi_awready  (sb_awready ),
      .sb_axi_awid     (sb_awid    ),
      .sb_axi_awaddr   (sb_awaddr  ),
      .sb_axi_awregion (sb_awregion),
      .sb_axi_awlen    (sb_awlen   ),
      .sb_axi_awsize   (sb_awsize  ),
      .sb_axi_awburst  (sb_awburst ),
      .sb_axi_awlock   (sb_awlock  ),
      .sb_axi_awcache  (sb_awcache ),
      .sb_axi_awprot   (sb_awprot  ),
      .sb_axi_awqos    (sb_awqos   ),
      .sb_axi_wvalid   (sb_wvalid  ),
      .sb_axi_wready   (sb_wready  ),
      .sb_axi_wdata    (sb_wdata   ),
      .sb_axi_wstrb    (sb_wstrb   ),
      .sb_axi_wlast    (sb_wlast   ),
      .sb_axi_bvalid   (sb_bvalid  ),
      .sb_axi_bready   (sb_bready  ),
      .sb_axi_bresp    (sb_bresp   ),
      .sb_axi_bid      (sb_bid     ),
      .sb_axi_arvalid  (sb_arvalid ),
      .sb_axi_arready  (sb_arready ),
      .sb_axi_arid     (sb_arid    ),
      .sb_axi_araddr   (sb_araddr  ),
      .sb_axi_arregion (sb_arregion),
      .sb_axi_arlen    (sb_arlen   ),
      .sb_axi_arsize   (sb_arsize  ),
      .sb_axi_arburst  (sb_arburst ),
      .sb_axi_arlock   (sb_arlock  ),
      .sb_axi_arcache  (sb_arcache ),
      .sb_axi_arprot   (sb_arprot  ),
      .sb_axi_arqos    (sb_arqos   ),
      .sb_axi_rvalid   (sb_rvalid  ),
      .sb_axi_rready   (sb_rready  ),
      .sb_axi_rid      (sb_rid     ),
      .sb_axi_rdata    (sb_rdata   ),
      .sb_axi_rresp    (sb_rresp   ),
      .sb_axi_rlast    (sb_rlast   ),

      //-------------------------- DMA AXI signals--------------------------
      .dma_axi_awvalid  (1'b0),
      .dma_axi_awready  (),
      .dma_axi_awid     (`RV_DMA_BUS_TAG'd0),
      .dma_axi_awaddr   (32'd0),
      .dma_axi_awsize   (3'd0),
      .dma_axi_awprot   (3'd0),
      .dma_axi_awlen    (8'd0),
      .dma_axi_awburst  (2'd0),

      .dma_axi_wvalid   (1'b0),
      .dma_axi_wready   (),
      .dma_axi_wdata    (64'd0),
      .dma_axi_wstrb    (8'd0),
      .dma_axi_wlast    (1'b0),

      .dma_axi_bvalid   (),
      .dma_axi_bready   (1'b0),
      .dma_axi_bresp    (),
      .dma_axi_bid      (),

      .dma_axi_arvalid  (1'b0),
      .dma_axi_arready  (),
      .dma_axi_arid     (`RV_DMA_BUS_TAG'd0),
      .dma_axi_araddr   (32'd0),
      .dma_axi_arsize   (3'd0),
      .dma_axi_arprot   (3'd0),
      .dma_axi_arlen    (8'd0),
      .dma_axi_arburst  (2'd0),

      .dma_axi_rvalid   (),
      .dma_axi_rready   (1'b0),
      .dma_axi_rid      (),
      .dma_axi_rdata    (),
      .dma_axi_rresp    (),
      .dma_axi_rlast    (),

      // clk ratio signals
      .lsu_bus_clk_en (1'b1),
      .ifu_bus_clk_en (1'b1),
      .dbg_bus_clk_en (1'b1),
      .dma_bus_clk_en (1'b1),

      .timer_int (timer_irq),
      .extintsrc_req ({4'd0, ethmac_irq, spi1_irq, spi0_irq, uart_irq}),

      .dec_tlu_perfcnt0 (),
      .dec_tlu_perfcnt1 (),
      .dec_tlu_perfcnt2 (),
      .dec_tlu_perfcnt3 (),

      .dmi_reg_rdata    (dmi_reg_rdata),
      .dmi_reg_wdata    (dmi_reg_wdata),
      .dmi_reg_addr     (dmi_reg_addr),
      .dmi_reg_en       (dmi_reg_en),
      .dmi_reg_wr_en    (dmi_reg_wr_en),
      .dmi_hard_reset   (dmi_hard_reset),

      .mpc_debug_halt_req (1'b0),
      .mpc_debug_run_req  (1'b0),
      .mpc_reset_run_req  (1'b1),
      .mpc_debug_halt_ack (),
      .mpc_debug_run_ack  (),
      .debug_brkpt_status (),

      .i_cpu_halt_req      (1'b0),
      .o_cpu_halt_ack      (),
      .o_cpu_halt_status   (),
      .o_debug_mode_status (),
      .i_cpu_run_req       (1'b0),
      .o_cpu_run_ack       (),

      .scan_mode  (1'b0),
      .mbist_mode (1'b0));

endmodule
