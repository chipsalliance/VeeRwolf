@00000000
0085051380001537
0285859300000597
0055002300058283
0005828300158593
800015B7FE029AE3
0005A02300958593
75462B5652657753
6F7220436F536573
000000000A736B63
