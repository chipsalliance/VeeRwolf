10008093030200B7
5041011307060137
908404130B0A1437
D0C484930F0E14B7
1FF0039300000193
0000023301000513
0021A2230011A023
0091A6230081A423
00028303004182B3
0012021302621C63
0001A023FEA218E3
0001A4230001A223
010181930001A623
80001537FC71C2E3
0010029301050513
0000006F00550023
0105051380001537
0055002300001337
000073B30012C293
FE731EE300138393
00000000FEDFF06F
