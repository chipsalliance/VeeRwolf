// SPDX-License-Identifier: Apache-2.0
// Copyright 2019 Western Digital Corporation or its affiliates.
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

//********************************************************************************
// $Id$
//
// Function: SweRVolf Nexys A7 clock generation
// Comments:
//
//********************************************************************************

module clk_gen_nexys
  (input      i_clk,
   input      i_rst,
   output     o_clk_core,
   output reg o_rst_core,
   output     o_clk50,
   output reg o_rst50
   );

   wire   clkfb;
   wire   locked;
   reg 	  locked_core_r;
   reg 	  locked50_r;

   wire   clock50_int;
   

   PLLE2_BASE
     #(.BANDWIDTH("OPTIMIZED"),
       .CLKFBOUT_MULT(16),
       .CLKIN1_PERIOD(10.0), //100MHz
       .CLKOUT0_DIVIDE(32),
       .CLKOUT1_DIVIDE(32),
       .DIVCLK_DIVIDE(1),
       .STARTUP_WAIT("FALSE"))
   PLLE2_BASE_inst
     (.CLKOUT0(o_clk_core),
      .CLKOUT1(clk50_int),
      .CLKOUT2(),
      .CLKOUT3(),
      .CLKOUT4(),
      .CLKOUT5(),
      .CLKFBOUT(clkfb),
      .LOCKED(locked),
      .CLKIN1(i_clk),
      .PWRDWN(1'b0),
      .RST(i_rst),
      .CLKFBIN(clkfb));

   BUFG BUFG_inst(.O(o_clk50),
		  .I(clk50_int)
		  );   

   always @(posedge o_clk_core) begin
      locked_core_r <= locked;
      o_rst_core <= !locked_core_r;
   end

   always @(posedge o_clk50) begin
      locked50_r <= locked;
      o_rst50  <= !locked50_r;
   end

endmodule
