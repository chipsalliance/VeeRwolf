0102829300000297
0600206F30529073
00112023FB010113
0041242300312223
0061282300512623
01C12C2300712A23
03E1202301D12E23
02A1242303F12223
02C1282302B12623
02E12C2302D12A23
0501202302F12E23
341022F305112223
300022F304512423
1BC000EF04512623
02051E6300000313
800003B7342022F3
0072F2B3FFF38393
00628A6300B00313
0000009700010513
78D0106F12408093
0042829304812283
0800006F04512423
0000639700010293
0043A1035D438393
00512023FF010113
001E0E130003AE03
3420257301C3A023
FFF28293800002B7
134000EF00557533
5902829300005297
00A282B300351513
0042A3030002A503
00006317000300E7
0003238358430313
00732023FFF38393
0002811300012283
02032E0300832383
00006297087E0863
0082A30355C28293
0293282302832623
03332C2303232A23
0553202303432E23
0573242305632223
0593282305832623
05B32C2305A32A23
0000639702232423
0003AE0309438393
0202A30307C32623
028321030062A423
0303248302C32403
0383298303432903
04032A8303C32A03
04832B8304432B03
05032C8304C32C03
05832D8305432D03
3412907304812283
3002907304C12283
0041218300012083
00C1228300812203
0141238301012303
01C12E8301812E03
02412F8302012F03
02C1258302812503
0341268303012603
03C1278303812703
0441288304012803
3020007305010113
00A312B300100313
000080673442B373
80000337342022F3
000005130062F2B3
0015051300028463
0000007300008067
4402829300006297
06C323830082A303
300522F300857513
0000806700038513
0200079302060063
00F04C6340C787B3
00000713FE060513
0007059300A5D533
00C5D73300008067
00F595B300C55533
FE9FF06F00B56533
0006081300058793
0005031300068713
000068B728069663
0EC5F6638B488893
0CE6786300010737
00C6B6B30FF00693
00D6573300369693
0008C70300E888B3
0200071300D706B3
00070C6340D70733
00D556B300E797B3
00F6E5B300E61833
0108551300E51333
0108161302A5F733
0103569301065613
0107171302A5D5B3
02B607B300D766B3
00F6FE6300058713
FFF58713010686B3
00F6F6630106E863
010686B3FFE58713
02A6F7B340F686B3
0103531301031313
0107979302A6D6B3
02D605B30067E333
00B37C6300068513
FFF6851300680333
00B3746301036663
01071713FFE68513
0000059300A76733
010007370E40006F
F2E66CE301000693
F31FF06F01800693
0010069300061663
000106B702C6D833
0FF006930CD87263
008007130106F463
00D888B300E856B3
00E686B30008C683
40D7073302000713
410787B30A071863
0108561300100593
0108D89301081893
02C7F73301035693
0107171302C7D7B3
02F8853300D766B3
00A6FE6300078713
FFF78713010686B3
00A6F6630106E863
010686B3FFE78713
02C6F7B340A686B3
0103531301031313
0107979302C6D6B3
02D888B30067E333
01137C6300068513
FFF6851300680333
0113746301036663
01071713FFE68513
0007051300A76733
010006B700008067
F4D862E301000713
F3DFF06F01800713
00D7D5B300E81833
00D556B300E51333
00E797B301085513
00F6E8B302A5F733
0107D79301081793
02A5D5B30108D613
00C7673301071713
0005861302B786B3
0107073300D77E63
01076863FFF58613
FFE5861300D77663
40D706B301070733
0108989302A6F733
02A6D6B30108D893
02D785B301071713
00068713011767B3
010787B300B7FE63
0107E863FFF68713
FFE6871300B7F663
40B787B3010787B3
00E5E5B301061593
18D5E663EB5FF06F
04E6F46300010737
00D835B30FF00813
0000673700359593
8B47071300B6D833
0007480301070733
0200059300B80833
02059663410585B3
EEF6ECE300100713
0016471300C53633
01000737EEDFF06F
FCE6E0E301000593
FB9FF06F01800593
00B696B301065733
0106DE9300D766B3
03D778B30107D733
0105583300B797B3
0106979300F86333
010358130107D793
03D7573300B61633
0108E83301089893
00070E1302E78F33
00D8083301E87E63
00D86863FFF70E13
FFE70E1301E87663
41E8083300D80833
03D8583303D878B3
03078EB301089893
0107D79301031793
0008071300F8E7B3
00D787B301D7FE63
00D7E863FFF80713
FFE8071301D7F663
010E1E1300D787B3
00010EB741D787B3
FFFE881300EE6733
0107589301077333
0106561301067833
0308883303030E33
02C30333010E5693
006686B301030333
0106F46302C888B3
0106D61301D888B3
0317E663011608B3
000107B7CF179AE3
00F6F6B3FFF78793
00FE7E3301069693
01C686B300B51533
DAD57CE300000593
CC9FF06FFFF70713
0000071300000593
FE010113DA5FF06F
00912A2300812C23
00112E2301212823
0005849300050913
56D030EF00060413
00A126231CD030EF
0010061300006537
BA45051300190593
00C12703458010EF
0000663706074263
BA060613000066B7
00006537BC868693
BB05051300090593
06040063430010EF
0487D6633E700793
F9C58593000065B7
0004851300040613
01812403410010EF
0141248301C12083
0000653701012903
02010113BF050513
000066373F00106F
B9C60613000066B7
FA1FF06FF9C68693
BC858593000065B7
000065B7FB9FF06F
00048513F9C58593
FB1FF06F3C0010EF
02912A23FC010113
02112E2303412423
0321282302812C23
0351222303312623
01712E2303612023
01912A2301812C23
01B1262301A12823
0005049300500793
0EF50E6300150A13
9B478793000067B7
00E7873300251713
002A171300072903
0007A98300E787B3
00006D3700006DB7
01900A9306400B13
00006C3700006CB7
0000061300006BB7
00048513B24D8593
FFF00593E95FF0EF
729010EF00090513
B3CD059300000613
E79FF0EF00048513
00098513FFF00593
529040EF70D010EF
B54C859303655433
0344043300048513
0014041301F47413
0004061303540433
00040513E45FF0EF
00098513379030EF
0000061318C020EF
00048513B6CC0593
00090513E25FF0EF
4D9040EF174020EF
B84B859303655433
0344043300048513
0014041301F47413
0004061303540433
00040513DF5FF0EF
F49FF06F329030EF
2909099300006937
2909091306498993
00006637F19FF06F
00006537000065B7
9CC60613FC010113
9DC505139D458593
02812C2302112E23
0321282302912A23
0341242303312623
0361202303512223
224010EF01712E23
0000643700001537
3885051300000593
44C020EF9B440413
0004250301840493
5F5010EF00440413
00006437FE941AE3
3084041300006937
000004936C090913
FFF00B9300300A93
0060099300400B13
0171222300000813
409A88B301612023
0004871300000793
300006137B000693
0004051300090593
001484935AD030EF
479030EF00040513
3009091307040413
03C12083FD3490E3
0341248303812403
02C1298303012903
02412A8302812A03
01C12B8302012B03
0000806704010113
0085530300452883
00A54F0300052803
FFF0079303130E33
0008859300F505A3
00C00F9300000613
01C8083302000E93
0000061301E64A63
0466CA6300000693
02BE57B300008067
03F6073300C52683
0047069300E68733
00D7242300D72223
00C505A300FEEC63
FFC5F5930025D593
FBDFF06F00160613
03D7C7B301F78793
0027979301072023
FDDFF06F00F80833
0005278300C52703
0047059300168693
00B7A02300C787B3
0116063300872583
0087258300B7A223
00F7242300F5A023
00058663F7DFF06F
0000806700C52223
0017F79300052783
00C5202300F66633
0005278300008067
00812C23FE010113
0121282300912A23
00112E2301312623
0005891300050993
0006041300F62023
0004258300100493
01C1208303259263
0004851301812403
0141248301012903
0201011300C12983
0049A78300008067
000780E700090513
00051E6300042783
004404130047A783
00148493FC0782E3
FB1FF06F00F42023
FFE7F7930007A783
00259793FE5FF06F
FF878793FD010113
00F50B3301612823
000B290303212023
0291222300478793
0281242300F504B3
0004A40300492783
0171262301412C23
0211262340F40A33
01512A2301312E23
08F41C63001A3B93
01403A3300442A83
0044298308F40C63
00B7DE6300200793
00040613FFCB2503
412585B300452583
ED1FF0EF0015B593
000B8593000A8613
EC1FF0EF00040513
000A059300090613
EB1FF0EF00040513
000B859300098613
EA1FF0EF00090513
008B202302C12083
0124A02302812403
0241248301C12983
01812A0302012903
01012B0301412A83
0301011300C12B83
00042A8300008067
F69FF06FFFEAFA93
FFE9F99300042983
0085A783F69FF06F
001787930005A703
00F5A42300279693
00A7202300D70733
001006930045A703
0007802300F707B3
0085A78300052503
FFE575130005A703
0027979300051A63
0007A50300F707B3
0017879300008067
00F5A42300279613
00A7202300C70733
00F707B30045A703
FBDFF06F00D78023
01712623FD010113
01312E2340000BB7
0181242301612823
0211262301A12023
0291222302812423
01412C2303212023
0191222301512A23
0005899300050D13
00100C1300060B13
0F3C5863FFFB8B93
002A1A1301798A33
FFCA2483014D0A33
0044AC83000A2903
001ABA9341990AB3
01991663000C8413
FFE474130004A403
0017F79300042783
0009859304079063
000D0513008A2023
0004A783DF5FF0EF
FFE7F79300198993
0004278300F4A023
0017E793000A2483
012A222300F42023
0044A40307990463
0044270300042A03
000A0863FFEA7A13
0017F793000A2783
0007086314078463
0017F79300072783
01691A6308078863
000A859300000613
CD9FF0EF00048513
FFE7F79300042783
0004A78300F42023
00070C630017F713
F29FF06FFFF98993
FFE474130004A403
0017E793F99FF06F
02C1208300F4A023
0241248302812403
01C1298302012903
01412A8301812A03
00C12B8301012B03
00412C8300812C03
0301011300012D03
0004278300008067
1080006FFFE7F793
0B990863000A0793
0007A68300070793
0A0692630016F693
000426830004A703
0017771300098593
00D76733FFE6F693
0004A70300E42023
00176713000D0513
0007A70300E4A023
00E7A02300176713
00FD07B300299793
CB1FF0EFFE87AE23
02812403F5691EE3
0201290302C12083
01812A0301C12983
00C12B8301012B03
00412C8300812C03
000A859300012D03
01412A8300048513
0000061302412483
BB9FF06F03010113
F79900E3000A0793
F4079CE300070793
00070A1301991463
FFCB8B9300299B93
008BA023017D0BB3
00198593014BA223
C31FF0EF000D0513
FFE7F79300042783
000A278300F42023
0017E793000BA403
EF990CE300FA2023
012BA02300442783
00052503F11FF06F
00058C6300050863
0007946300452783
0007851300008067
00052783FE9FF06F
FE9FF06FFFE7F793
02812423FD010113
01312E2302912223
0321202302112623
01512A2301412C23
0171262301612823
0005A78303010413
000509930005A223
00F5A0230017F793
0005849300052783
00B9A02304079263
00F5242300100793
FD04011300F5A023
0281240302C12083
0201290302412483
01812A0301C12983
01012B0301412A83
0301011300C12B83
0085278300008067
0027979300010A93
FF07F79301378793
00010A1340F10133
A99FF0EF000A0613
00FA093300251793
0049A783FFC92B83
000B859300050B13
000780E700048513
0004861300154593
0FF5F593000B8513
0004A783A45FF0EF
00992023001B0B13
00F4A023FFE7F793
00090793000B0B93
01784A6300100813
00072783000A2703
0CC0006F0017E793
FFC78913FFC7A603
0017771300062703
FF87A5830A071E63
0045A703FF878493
00E6166300070693
FFE6F6930005A683
0006A50304068063
0015751300048793
0005A70302051863
FFE77713FFEB8B93
0006270300E5A023
00E6202300176713
001767130006A703
F81FF06F00E6A023
00FA07B3002B9793
00462683FFC7A783
0017371340E60733
0017B79340D787B3
000B859300F70863
A21FF0EF000A0513
000A0513FFFB8593
0004A703A15FF0EF
0017E79300072783
0009270300F72023
FFE7F79300072783
0089A78300F72023
0169A4230167D463
00F9A023000A2783
E61FF06F000A8113
02812423FD010113
01412C2302912223
0171262301612823
0211262301812423
01312E2303212023
0191222301512A23
0085278303010413
00050B1300010B93
0137879300279793
40F10133FF07F793
000A061300010A13
8E9FF0EF00058493
018A0C3300251C13
10979263FFCC2783
000509930004A903
0C090463FFE97913
0C0780630044A783
0000051300100793
FF8C25030137D463
00198713012C2023
00271A9300492783
015A0AB300070993
FF8AAC830E079E63
0045258310050263
409585B300090613
859FF0EF0015B593
000927030F949A63
FFE777130004A783
00E7E7B30017F793
0009278300F4A023
00F4E7B30017F793
0044A78300F92023
FFCAA70300F92223
0004A223FFCC2783
FEFAAE23FEEC2E23
000927030004A683
00177713FFE6F793
00E4A02300F76733
0016F69300092783
00D7E7B3FFE7F793
0004A78300F92023
00091463FFE7F913
001007130044A903
012B20230B374C63
000927830A090463
00F920230017E793
FD040113000B8113
0281240302C12083
0201290302412483
01812A0301C12983
01012B0301412A83
00812C0300C12B83
0301011300412C83
00FAA02300008067
0007891300170713
012B2023EE9FF06F
004CA583F11FF06F
000C851300048613
0015B593412585B3
0004A703F4CFF0EF
0017779300092683
00D7E7B3FFE6F693
0009278300F4A023
0017F793FFE77713
EF5FF06F00E7E7B3
F65FF06F000B2423
015A0AB300299A93
02091863FF8AA503
000486130017F793
0045258306079463
409585B300000613
EE8FF0EF0015B593
00FB2023000A2783
00452583F29FF06F
409585B300090613
EC8FF0EF0015B593
0017F7930004A783
0009278300078863
00079A630017F793
0017E79300092783
FBDFF06F00F92023
00000613FF2AAE23
000A051300098593
FA5FF06F8B1FF0EF
0005879300052503
0000051300051663
0085A68300008067
00E69463FFF00713
0005A603815FF06F
00E6073300269713
0045250300072503
0045A583FE0514E3
0005450300D58533
FFF6869300050C63
FFC7250300D7A423
00E7A42300008067
FFF687130087A683
00D586B300D05863
FE0684E30006C683
F80748E300E7A423
00E6073300271713
0000806700072503
00050793FF010113
0006059300058513
0011262300068613
76D020EF000780E7
00000513620030EF
FF01011300008067
0005041300812423
0011262304500513
0005849300912223
00048593000400E7
000400E705200513
0081240300040313
0004859300C12083
0520051300412483
0003006701010113
001787930005A783
000067B700F5A023
000300671F07A303
04812423FB010113
03412C2303312E23
0371262303512A23
0491222304112623
0361282305212023
0391222303812423
01B12E2303A12023
00058A9300050A13
00068B9300060993
00E0546300100413
0010079300070413
00FB946302000C13
3B9AD4B703000C13
00A00B1300100913
A004849300000793
00200D9300100C93
0007946300A00D13
0299D5330899E063
00190913000A8593
000A00E703050513
FFFB0B1300100793
03A4D4B30299F9B3
000A8593FD9B1AE3
000A00E703098513
4124043300300793
04C1208306FB8A63
0441248304812403
03C1298304012903
03412A8303812A03
02C12B8303012B03
02412C8302812C03
01C12D8302012D03
0000806705010113
F97DECE3F9644EE3
000C0513000A8593
000A00E700F12623
00C1278300190913
000A8593F7DFF06F
000A00E702000513
FE8048E3FFF40413
000067B7F8DFF06F
000080671EA7A823
04812423FB010113
0521202304912223
03412C2303312E23
03A1202303512A23
0411262301B12E23
0371262303612823
0391222303812423
0005849300050413
00068D9300060A93
FFF0099300000913
00000D1300000A13
04051063000AC503
0481240304C12083
0401290304412483
03812A0303C12983
03012B0303412A83
02812C0302C12B83
02012D0302412C83
0501011301C12D83
000D1E6300008067
3AD5086302500693
000400E700048593
FA5FF06F001A8A93
12D50E6306400693
0390069306A6E263
0310069302A6EA63
02D006930ED57C63
0300079338D50863
025007130CF50863
0004859302E51263
000400E702500513
0580069318C0006F
063007131ED50663
0004859332E50A63
000400E702500513
000AC50300048593
07000693FD5FF06F
02A6E8631AD50263
0CD5026306900693
00D5066306C00693
FCD514E306800693
08D51A6306800693
0480091308A91E63
07500693F59FF06F
02A6EE6312D50663
FAE510E307300713
004D8B93000DAC03
000B4503000C0B13
0030079328051C63
418B0B3300FA1863
29604A6341698B33
0E80006F000B8D93
14D5046307800693
F99FF06F07A00693
2A0A0E630009DE63
EE0A1AE3FD050993
EEDFF06F00200A13
00A00693FE09C8E3
FD09899302D989B3
FE1FF06F013509B3
00D5146306C00693
F20910E328A90863
EBDFF06F00050913
04E9126307A00713
004D8D93000DA603
0004859302065063
00C1242302D00513
00812603000400E7
40C00633FFF98993
000A069300098713
0004051300048593
0480006FC79FF0EF
FAE90EE306C00713
FAE91AE304C00713
FF87F713007D8793
0047268300072603
8000073700870D93
00C7373300E60733
F8070AE300D70733
0004051300048593
00000D13BCDFF0EF
07A00713E29FF06F
000DA60300E91863
F8DFF06F004D8D93
FEE908E306C00713
FEE914E304C00713
FF87F713007D8793
0007260300870D93
F60702E300472703
00048593FB1FF06F
000400E703000513
0780051300048593
00800993000400E7
000AC60300100A13
00D61A6307000693
00000C13000DAB83
0280006F004D8D93
FED906E306C00693
FED912E304C00693
FF87F693007D8793
0046AC030006AB83
0100079300868D93
0001242300000C93
FFCB0B1304000B13
000B8513000B0613
00F12623000C0593
00F57513861FE0EF
0605166300C12783
0300069300812703
060B186300071463
0185151300A68533
4185551300048593
000400E700F12423
00812783001C8C93
00300693020B1863
D0DA1AE300000D13
41970CB300199713
00048593ED905EE3
000400E702000513
FEDFF06FFFFC8C93
F79FF06F01A12423
0570069300900713
03000693FAA760E3
FFF78713F99FF06F
00F9CC6300E12623
00FA1C6300100793
0300051300048593
00C12783000400E7
00200793F3DFF06F
00048593FEFA1AE3
FE5FF06F02000513
001B0B1300048593
D59FF06F000400E7
0200051300048593
FFFB0B13000400E7
000DA503D5DFF06F
00048593004D8B13
000B0D93000400E7
00000913E35FF06F
00000A13FFF00993
C4DFF06F00100D13
C45FF06F00300A13
C3DFF06F00100A13
C35FF06F04C00913
00050613FE010113
0005869300001537
00C1059355050513
0001262300112E23
01C12083B61FF0EF
0000806702010113
02B12223FC010113
00112E2302410593
02D1262302C12423
02F12A2302E12823
03112E2303012C23
FA5FF0EF00B12623
0401011301C12083
000065B700008067
FF01011300006537
BE850513BCC58593
0011262302700613
00C12083FA9FF0EF
0040051300000593
1090006F01010113
0080079300008067
304050733007B7F3
0000806734405073
00812423FF010113
0000643700912223
00A0079300112623
2684041300050493
0004250300F51C63
00D0059300452783
000780E70047A783
0045278300042503
0047A7830FF4F593
00C12083000780E7
0004851300812403
0101011300412483
0000253700008067
A51FF06FBF050513
00112623FF010113
BF45051300006537
000067B77B8000EF
FD9FF0EF26A7A423
0000051300C12083
0000806701010113
0007A023F00C37B7
00478713F00C27B7
0007202312C78793
FEF71CE300470713
00478713F00C07B7
12C7879300F00693
0047071300D72023
F00C47B7FEF71CE3
12C7879300478713
0047071300072023
F00C57B7FEF71CE3
12C7879300478713
0047071300072023
BC905073FEF71CE3
BCC05073BCB05073
80078793000017B7
000005133047A7F3
FF01011300008067
0081242300112623
FC802473BCA05073
0FF4741300245413
2687A623000067B7
03E00793FFF40713
0000051300E7F663
00B407132F0000EF
00371713000057B7
00E787B367878793
000706630047A703
000700E70007A503
40B78793000017B7
0024141300F40433
00F40433F00C07B7
00C1208300042023
0101011300812403
FF55071300008067
02E7E66303F00793
3007B7F300800793
F00C07377F550513
00E5053300251513
00E5202300100713
3007A7F30087F793
00B0071300008067
00A7746300050793
00100513FBDFF06F
3045257300F51533
800017B700008067
0207A5030247A703
FEE59AE30247A583
FE01011300008067
00112E2300912A23
0121282300812C23
0141242301312623
0161202301512223
3004B4F300800493
2709051300006937
784020EF0084F493
0000643702051E63
00006537000065B7
04F00693C2458593
C3C50513C0840613
00006537CF9FF0EF
CEDFF0EFC5C50513
C084051304F00593
27090513D1DFF0EF
794020EF00006AB7
F61FF0EF258A8A93
004AAB03000AA403
4085053300050A13
0005899300AA37B3
416585B30007A637
0000069312060613
BD4FE0EF40F585B3
120787930007A7B7
0085073302F50533
00A7353300F707B3
00E7B633016506B3
41478A3300D60633
413609B30147B5B3
00DAA22300EAA023
0330426340B989B3
3E70059300099663
000F47B70145EC63
00F707B324078793
00D7063300E7B733
FFF0069380001737
02F7242302D72623
2709051302C72623
02051E636B0020EF
000065B700006437
C745859300006537
C084061306200693
BFDFF0EFC3C50513
C8C5051300006537
06200593BF1FF0EF
C21FF0EFC0840513
018124033004A4F3
0141248301C12083
00C1298301012903
00412A8300812A03
0010051300012B03
2740306F02010113
00112623FF010113
0007A7B7E3DFF0EF
8000173712078793
FFF0069300F507B3
00A7B53302D72623
02F7242300B50533
0070051302A72623
00C12083DEDFF0EF
0101011300000513
0000806700008067
0000806700000513
3007A7F300800793
FF01011300008067
4B8000EF00112623
00112623FF010113
342027F300050593
4A0000EF00000513
00112623FF010113
00000593342027F3
FC9FF0EF00100513
00112623FF010113
B79FF0EF530000EF
F14025735A4000EF
1050007300050663
00006117FFDFF06F
000012B7E4410113
0051013380028293
C44FF06FFC9FF0EF
02812423FD010113
0321202302912223
01412C2301312E23
0161282301512A23
0211262301712623
0181242300078B93
0005099302800793
0006049300058413
00070B1300068A13
0008891300080A93
000027B708F89863
08F6986356078793
0004059303012703
0004861300090693
380020EF00098513
00B405B3FB048593
FF05F593000027B7
04F5A62388078793
02C12083000027B7
0947879302812403
0365A6230345A423
0355AA230375A823
02B9A42304F5A423
0201290302412483
01812A0301C12983
01012B0301412A83
00812C0300C12B83
0000806703010113
0440079301D88713
00006C37F6E7FCE3
00006537000065B7
01500693CA0C0613
C3C50513CC858593
000065379C9FF0EF
FE30069300090593
D5C5051302700613
015005939B1FF0EF
9E1FF0EFCA0C0513
00054783F31FF06F
00E794630005C703
40E7853300079663
0015051300008067
FE1FF06F00158593
000507930FF5F693
040718630037F713
008597130FF5F593
0105971300B765B3
00C7833300B765B3
0030081300078713
03186E6340E308B3
0027159300265713
FFC0059300B787B3
00C7073302B70733
02E7946300E78733
FE060EE300008067
FED78FA300178793
F9DFF06FFFF60613
FEB72E2300470713
00178793FB9FF06F
FD1FF06FFED78FA3
0080071300852803
0048268330073773
0606886300877713
0087A78300052783
060600630007A603
00C787B300369793
0085288302D7D7B3
00C5C6030008A583
080663130FF67613
0085230300658623
0047D59300032303
00B300230FF5F593
00C7D79300852583
0005A5830FF7F793
0085278300F58223
00C786230007A783
0085278300D8A223
0007A78300300693
0088478300D78623
0017F79300B00693
02B0069300078463
0007A78300852783
0085278300D78823
0007A783F8700693
0085278300D78423
0007C6830007A783
3007277300078223
0000806700000513
0007A70300852783
0017F79301474783
0007478300078A63
00F5802300000513
FFF0051300008067
0085278300008067
014706930007A703
0207F7930006C783
00B70023FE078CE3
0085278300008067
0147C5030007A783
00F5751300155513
0025171300008067
00150513000067B7
00251513DA478793
00E78733FF010113
0081242300A787B3
0007240300912223
001126230007A483
00C1208300946C63
0041248300812403
0000806701010113
0004051300042783
000780E70047A783
0004222300050463
FCDFF06F00C40413
000067B7FF010113
000064B700912223
0011262300812423
0121202320478413
2404849320478793
0005091300941C63
0294146300078413
0440006F00000413
0007086300442703
0007270300042703
00C4041302A70863
00442783FD1FF06F
00C4041300079663
00042783FCDFF06F
0007A58300090513
FE0514E3D2DFF0EF
00C1208300040513
0041248300812403
0101011300012903
0080079300008067
0000006F3007B7F3
00112623FF010113
FE010113FEDFF0EF
00112E2300812C23
0005041300912A23
76D010EF00B12623
0005049300C12583
FCDFF0EF00040513
02F41E6300400793
000065B700006437
DD45859300006537
DB84061308700693
E3CFF0EFC3C50513
DF45051300006537
08700593E30FF0EF
E60FF0EFDB840513
01C1208301812403
0141248300048513
5BC0206F02010113
00812423FF010113
0080041300112623
2D5020EF300437F3
0010051300A04463
3A1020EF00100593
FE5FF06FA89FF0EF
000067B700006537
6BC7879325850613
0000059340C78633
C45FF06F25850513
00200513FF010113
E01FF0EF00112623
000065B700006637
F9C6061300006537
E4C50513E2C58593
00300513D90FF0EF
2A0020EFDDDFF0EF
000067B7B1CFE0EF
00C7C70361878793
00E78623FFE77713
0101011300C12083
F601011300008067
000087B708812C23
0931262300006437
688409936C078793
0101079300F9A223
0000059307000613
08112E2300078513
0921282308912A23
BA5FF0EF09412423
00A9A42300100A13
01410EA300000513
00100513D5DFF0EF
10100793D55FF0EF
225010EF00F11E23
00006937000067B7
000026B7E7478793
61890493000085B7
0000071300F12223
0141202300000793
0000081300000893
400006135B068693
618905138C058593
5F9010EF0299A023
6884041300D4C783
00E486A3FFB7F713
00079A6301B7F793
000796630184A783
170010EF61890513
E7C78793000067B7
0000653700F12223
000026B700100793
5A850493000085B7
0280089300F12023
0000079300000813
5606869300000713
CC05859320000613
589010EF5A850513
0094262300D4C783
FFB7F79300800513
000067B700F486A3
00F42C236A078793
3005357300F42E23
AE9FD0EF00857513
0005262300052423
00A5222300A52023
FE01011300008067
0121282300912A23
00112E2301412423
0131262300812C23
00058A1300050493
3009397300800913
2744051300006437
625010EF00897913
000069B702051E63
00006537000065B7
04F00693C2458593
C3C50513C0898613
00006537B98FF0EF
B8CFF0EFC5C50513
C089851304F00593
27440513BBCFF0EF
00C4A703639010EF
68878793000067B7
0084A50306070263
0ED500630087A683
274405130E0A1263
02051E635E1010EF
000065B700006437
C745859300006537
C084061306200693
B2CFF0EFC3C50513
C8C5051300006537
06200593B20FF0EF
B50FF0EFC0840513
FF00051330092973
0087A68306C0006F
0087A78300E68683
00D4A82300170713
00F4A42300E4A623
575010EF27440513
0000643702051E63
00006537000065B7
06200693C7458593
C3C50513C0840613
00006537AC0FF0EF
AB4FF0EFC8C50513
C084051306200593
30092973AE4FF0EF
01C1208300000513
0141248301812403
00C1298301012903
0201011300812A03
0104A68300008067
00E50783F7DFF06F
00B7D46300E68583
0005D46300078593
0000099300000593
644010EF00F5D663
000A069300050993
0009059300048613
5A4010EF27440513
00800913F8050EE3
2744051330093973
48D010EF00897913
00006A3702051E63
00006537000065B7
04F00693C2458593
C3C50513C08A0613
00006537A00FF0EF
9F4FF0EFC5C50513
C08A051304F00593
27440513A24FF0EF
0004A7834A1010EF
00F48E630104A583
00E7878300078C63
0007859300B7D463
000005930005D463
00E507830084A503
0209826300F59E63
2744051300090593
FF5005135EC000EF
584010EFEFDFF06F
FE1FF06FFE0514E3
415010EF27440513
0000643702051E63
00006537000065B7
06200693C7458593
C3C50513C0840613
00006537960FF0EF
954FF0EFC8C50513
C084051306200593
30092973984FF0EF
00C52783FA5FF06F
00812C23FE010113
00912A2300112E23
0131262301212823
02079E6300050413
000065B7000064B7
EA05859300006537
E84486130D300693
8FCFF0EFC3C50513
EB85051300006537
0D3005938F0FF0EF
920FF0EFE8448513
68848793000064B7
0087A78300842703
02F70E6368848493
000065B700006937
EBC5859300006537
E84906130D400693
8ACFF0EFC3C50513
EB85051300006537
0D4005938A0FF0EF
8D0FF0EFE8490513
02078E630004A783
000065B700006937
F005859300006537
EDC9061310C00693
86CFF0EFC3C50513
EB85051300006537
10C00593860FF0EF
890FF0EFEDC90513
00F7C7030084A783
02F71E6300100793
000065B700006937
F145859300006537
EDC9061310D00693
824FF0EFC3C50513
EB85051300006537
10D00593818FF0EF
848FF0EFEDC90513
00F747830084A703
00F707A3FFF78793
0010071300C42783
FFF7879302E78463
0181240300F42623
0141248301C12083
00C1298301012903
3390006F02010113
3004B4F300800493
2749051300006937
21D010EF0084F493
000069B702051E63
00006537000065B7
04F00693C2458593
C3C50513C0898613
00006537F91FE0EF
F85FE0EFC5C50513
C089851304F00593
27490513FB5FE0EF
00842503231010EF
00E5078301042583
34C010EF00F58463
6B4000EF00040513
02050C6300A42423
00E4282300E50703
0605262300D54703
0007186301F77713
0007946301852783
00048593415000EF
368000EF27490513
00042623F35FF06F
19D010EF27490513
0000643702051E63
00006537000065B7
06200693C7458593
C3C50513C0840613
00006537EE9FE0EF
EDDFE0EFC8C50513
C084051306200593
3004A4F3F0DFE0EF
00D54783EE5FF06F
0007986301F7F793
0015351301852503
0000051300008067
00E5070300008067
0010079300E58683
0000079300D74C63
0105278300E6C863
00A7B7B30105A503
0000806700078513
FF01011300052783
0011262300812423
0005041300912223
000064B702079863
00006537000065B7
C3C50513FBC58593
FA0486131AE00693
1AE00593E41FE0EF
E71FE0EFFA048513
00C1208300042503
0041248300812403
0000806701010113
00812423FF010113
2804041300006437
0011262300042783
A9CFF0EF02078863
0081240300042783
00A7853300C12083
68A72C2300006737
0007851300000593
3900206F01010113
0081240300C12083
0000806701010113
00812C23FE010113
0141242301212823
00912A2300112E23
0005091301312623
0080041300058A13
000064B730043473
0084741327848513
02051E637F0010EF
000065B7000069B7
C245859300006537
C089861304F00693
D65FE0EFC3C50513
C5C5051300006537
04F00593D59FE0EF
D89FE0EFC0898513
005010EF27848513
6807AC23000067B7
00A0079300990913
000067B702F95933
000067B72927A023
F05FF0EF2747AE23
7A4010EF27848513
000064B702051E63
00006537000065B7
06200693C7458593
C3C50513C0848613
00006537CF1FE0EF
CE5FE0EFC8C50513
C084851306200593
30042473D15FE0EF
0181240301C12083
0101290301412483
00812A0300C12983
0000806702010113
00812C23FE010113
00112E2301212823
0131262300912A23
0080041300050913
000064B730043473
0084741327848513
02051E636E8010EF
000065B7000069B7
C245859300006537
C089861304F00693
C5DFE0EFC3C50513
C5C5051300006537
04F00593C51FE0EF
C81FE0EFC0898513
6FC010EF27848513
DBDFF0EF00890513
300000EF00090593
2784851300D94783
00F906A3FFD7F793
02051E636A8010EF
000065B7000064B7
C745859300006537
C084861306200693
BF5FE0EFC3C50513
C8C5051300006537
06200593BE9FE0EF
C19FE0EFC0848513
01C1208330042473
0009242301812403
0101290301412483
0201011300C12983
FF01011300008067
0011262300812423
0085F41300912223
0604066300050793
6887270300006737
0005849306071063
02051E63618010EF
000065B700006437
C745859300006537
C084061307900693
B65FE0EFC3C50513
C8C5051300006537
07900593B59FE0EF
B89FE0EFC0840513
00C1208300812403
0041248300048513
A10FD06F01010113
5BC010EF00078513
000064B702051E63
00006537000065B7
06200693C7458593
C3C50513C0848613
00006537B09FE0EF
AFDFE0EFC8C50513
C084851306200593
30042473B2DFE0EF
0081240300C12083
0101011300412483
0085779300008067
0000673700078A63
0007146368872703
3007A7F399CFD06F
0080051300008067
0085751330053573
FE010113FD5FF06F
00112E2300812C23
0121282300912A23
0080041301312623
000064B730043473
0084741327848513
02051E634E0010EF
000065B700006937
C245859300006537
C089061304F00693
A55FE0EFC3C50513
C5C5051300006537
04F00593A49FE0EF
A79FE0EFC0890513
0000693727848513
688927834F0010EF
02078E6368890913
000065B7000069B7
F005859300006537
EDC9861310C00693
A05FE0EFC3C50513
EB85051300006537
10C005939F9FE0EF
A29FE0EFEDC98513
00F7C70300892783
02F71E6300100793
000065B7000069B7
F145859300006537
EDC9861310D00693
9BDFE0EFC3C50513
EB85051300006537
10D005939B1FE0EF
9E1FE0EFEDC98513
00F7478300892703
00F707A3FFF78793
41C010EF27848513
000064B702051E63
00006537000065B7
06200693C7458593
C3C50513C0848613
00006537969FE0EF
95DFE0EFC8C50513
C084851306200593
3004247398DFE0EF
0181240301C12083
0101290301412483
0201011300C12983
FF01011300008067
00812423000067B7
0091222300112623
000584135A878793
000064B702F59863
00006537000065B7
C3C50513FF458593
FA0486132C100693
2C1005938F1FE0EF
921FE0EFFA048513
0004278300442703
0041248300C12083
00E7A22300F72023
0004222300042023
0101011300812403
0005278300008067
0000079300F51463
0000806700078513
01212823FE010113
00112E2301312623
00912A2300812C23
0080091300050993
000064B730093973
0089791327848513
02051E632D8010EF
000065B700006437
C245859300006537
C084061304F00693
84DFE0EFC3C50513
C5C5051300006537
04F00593841FE0EF
871FE0EFC0840513
2EC010EF27848513
F71FF0EF00098513
2784851300050413
02051E632A8010EF
000065B7000069B7
C745859300006537
C089861306200693
FF4FE0EFC3C50513
C8C5051300006537
06200593FE8FE0EF
819FE0EFC0898513
0C04066330092973
3009397300800913
0089791327848513
02051E63228010EF
000065B7000069B7
C245859300006537
C089861304F00693
F9CFE0EFC3C50513
C5C5051300006537
04F00593F90FE0EF
FC0FE0EFC0898513
23C010EF27848513
8FDFF0EF00840513
E41FF0EF00040593
2784851300D44783
00F406A3FFD7F793
02051E631E8010EF
000065B7000064B7
C745859300006537
C084861306200693
F34FE0EFC3C50513
C8C5051300006537
06200593F28FE0EF
F58FE0EFC0848513
0004242330092973
2F5010EF01840513
01C1208300040513
0141248301812403
00C1298301012903
0000806702010113
02812423FD010113
0321202302912223
01312E2302112623
000067B703010413
000504935A878793
02F5986300058913
000065B7000069B7
FF45859300006537
2E500693C3C50513
E9CFE0EFFA098613
FA0985132E500593
00C4A703ECCFE0EF
00F4A62300170793
04079A6300E92823
002797130084A783
FF07771301770713
40E1013301778793
00F10713FF07F793
00F1079340F10133
FF077713FF07F793
FFF00793FCF42C23
FCF42E23FCE42A23
00048513FD440593
02051863F11FD0EF
0004851300090593
FD040113A61FD0EF
0281240302C12083
0201290302412483
0301011301C12983
00C4A78300008067
00E4A62300178713
FB5FF06F00F52823
000067B7FF010113
0091222300812423
0121202300112623
000504135A878793
02F5986300058493
000065B700006937
FF45859300006537
30000693C3C50513
DA4FE0EFFA090613
FA09051330000593
00048593DD4FE0EF
BCDFD0EF00040513
0007946300042783
00C1208300042623
0041248300812403
0101011300012903
0000059300008067
FF010113975FD06F
0000643700812423
0005091301212023
0245051368840513
0011262300912223
68840413FD5FF0EF
0005146300050493
06091E6300C42483
02079E6300842783
000065B700006937
FD45859300006537
FA09061307500693
CFCFE0EFC3C50513
EB85051300006537
07500593CF0FE0EF
D20FE0EFFA090513
00D7C70300842783
0207166301F77713
07F0071300E7D683
02F4202302D77063
0081240300C12083
0001290300412483
0000806701010113
0097846300842783
02942023E88FF0EF
FE010113FD9FF06F
0000693701212823
0087A78368890793
00812C2300112E23
00912A2300F7C783
6889091301312623
0000643702079E63
00006537000065B7
25800693F3C58593
C3C50513FA040613
00006537C48FE0EF
C3CFE0EFEB850513
FA04051325800593
00092783C6CFE0EF
0000643702078E63
00006537000065B7
25900693F0058593
C3C50513FA040613
00006537C08FE0EF
BFCFE0EFEB850513
FA04051325900593
00800413C2CFE0EF
000064B730043473
0084741327848513
02051E63641000EF
000065B7000069B7
C245859300006537
C089861304F00693
BB4FE0EFC3C50513
C5C5051300006537
04F00593BA8FE0EF
BD8FE0EFC0898513
655000EF27848513
0000051300892703
0017879300F74783
E21FF0EF00F707A3
605000EF27848513
000064B702051E63
00006537000065B7
06200693C7458593
C3C50513C0848613
00006537B50FE0EF
B44FE0EFC8C50513
C084851306200593
30042473B74FE0EF
01C1208301812403
0101290301412483
0201011300C12983
FE010113865FF06F
0121282300812C23
00912A2300112E23
0005091301312623
3004347300800413
27848513000064B7
54D000EF00847413
000069B702051E63
00006537000065B7
04F00693C2458593
C3C50513C0898613
00006537AC0FE0EF
AB4FE0EFC5C50513
C089851304F00593
27848513AE4FE0EF
00006537561000EF
6AC5051300090593
00D94783BA9FF0EF
0407E79300000513
D21FF0EF00F906A3
505000EF27848513
000064B702051E63
00006537000065B7
06200693C7458593
C3C50513C0848613
00006537A50FE0EF
A44FE0EFC8C50513
C084851306200593
30042473A74FE0EF
0181240301C12083
0101290301412483
0201011300C12983
FF05278300008067
00812C23FE010113
00112E2301312623
0121282300912A23
0005041301412423
0C078463FE850993
3004B4F300800493
2789051300006937
43D000EF0084F493
00006A3702051E63
00006537000065B7
04F00693C2458593
C3C50513C08A0613
000065379B0FE0EF
9A4FE0EFC5C50513
C08A051304F00593
278905139D4FE0EF
FF040513451000EF
00098593B10FF0EF
FF544783855FF0EF
FFD7F79327890513
3FD000EFFEF40AA3
0000693702051E63
00006537000065B7
06200693C7458593
C3C50513C0890613
00006537948FE0EF
93CFE0EFC8C50513
C089051306200593
3004A4F396CFE0EF
FF544783FE042823
FEB7F79300098513
A50FF0EFFEF40AA3
0181240302050463
0141248301C12083
00812A0301012903
00C1298300098513
DD9FF06F02010113
0181240301C12083
0101290301412483
00812A0300C12983
0000806702010113
00812C23FE010113
00112E2301212823
0131262300912A23
0080041300050913
000064B730043473
0084741327848513
02051E63301000EF
000065B7000069B7
C245859300006537
C089861304F00693
874FE0EFC3C50513
C5C5051300006537
04F00593868FE0EF
898FE0EFC0898513
315000EF27848513
0000653700D94783
0407F7936AC50993
0009059300078863
A4DFF0EF6AC50513
0009851300090593
00D94783941FF0EF
00F906A30407E793
68878793000067B7
412505330087A503
AA9FF0EF00153513
28D000EF27848513
000064B702051E63
00006537000065B7
06200693C7458593
C3C50513C0848613
00006537FD9FD0EF
FCDFD0EFC8C50513
C084851306200593
30042473FFDFD0EF
0181240301C12083
0101290301412483
0201011300C12983
000067B700008067
000067B72807A703
0607046368878793
07F006930087A703
04C6EC6300E75603
00E70603000066B7
04D6446327C6A683
5A86061300006637
0187268302C70E63
0107A68302069A63
FF01011302D54063
0011262300070513
00C12083E79FF0EF
91CFF06F01010113
00D7A82340A686B3
0007A82300008067
FE01011300008067
0131262300812C23
00912A2300112E23
0005099301212823
3004347300800413
27848513000064B7
155000EF00847413
0000693702051E63
00006537000065B7
04F00693C2458593
C3C50513C0890613
00006537EC9FD0EF
EBDFD0EFC5C50513
C089051304F00593
27848513EEDFD0EF
00D9C783169000EF
6889091300006937
00078E630407F793
0249051300098593
00D9C7838A1FF0EF
00F986A3FBF7F793
4135053300892503
911FF0EF00153513
0F5000EF27848513
000064B702051E63
00006537000065B7
06200693C7458593
C3C50513C0848613
00006537E41FD0EF
E35FD0EFC8C50513
C084851306200593
30042473E65FD0EF
0181240301C12083
0101290301412483
0201011300C12983
FE01011300008067
00912A2300812C23
0121282300050413
0131262300112E23
0006049300058913
00D44783EC5FF0EF
00F406A30027E793
000067B706090663
5A87879301242423
000069B702F41863
00006537000065B7
C3C50513FF458593
FA0986132AB00693
2AB00593DA1FD0EF
DD1FD0EFFA098513
0AF90E6300092783
00E407030A078C63
08D75E6300E78683
00F420230047A703
0087202300E42223
FFF007930087A223
0204DE630AF48663
000065B700006937
F645859300006537
FA09061319800693
D3DFD0EFC3C50513
F745051300006537
19800593D31FD0EF
D61FD0EFFA090513
000004930004D463
00A0061300948493
0184051302C4D633
01C1208301812403
0101290301412483
000045B700C12983
0201011395458593
6A10006F00160613
00D7866300492683
F4079AE30007A783
0124202300492783
0049278300F42223
008922230087A023
01C12083F55FF06F
0141248301812403
00C1298301012903
0000806702010113
000067B7FF010113
0005041300812423
009122236907A503
0006059300058493
0011262300068613
00040513E6DFF0EF
02051E636F8000EF
000065B700006437
C745859300006537
C084061307900693
C45FD0EFC3C50513
C8C5051300006537
07900593C39FD0EF
C69FD0EFC0840513
00C1208300812403
0041248300048513
AF0FC06F01010113
00812C23FE010113
0131262301212823
00912A2300112E23
0151222301412423
0005899300050913
3004347300800413
27848513000064B7
63C000EF00847413
00006A3702051E63
00006537000065B7
04F00693C2458593
C3C50513C08A0613
00006537BB1FD0EF
BA5FD0EFC5C50513
C08A051304F00593
27848513BD5FD0EF
00090513650000EF
01899993CC5FE0EF
4189D99300050A93
00006A370A050063
000905936ACA0A13
D7CFF0EF000A0513
01390723000A0513
C6CFF0EF00090593
DF0FF0EF00100513
5D4000EF27848513
000064B702051E63
00006537000065B7
06200693C7458593
C3C50513C0848613
00006537B21FD0EF
B15FD0EFC8C50513
C084851306200593
30042473B45FD0EF
0181240301C12083
01412483000A8513
00C1298301012903
00412A8300812A03
0000806702010113
F8DFF06F01390723
00003737000067B7
CC47071368878793
0000051300000593
0207A6230207A223
02E7A4230207A823
00E50503CE9FE06F
FE01011300008067
0000643700812C23
00112E2368842783
0121282300912A23
6884041301312623
000064B702078E63
00006537000065B7
3B500693F0058593
C3C50513FA048613
00006537A59FD0EF
A4DFD0EFEB850513
FA0485133B500593
00842703A7DFD0EF
5A878793000067B7
008007930CF70E63
000064B73007B7F3
0087F99327848513
02051E63480000EF
000065B700006937
C245859300006537
C089061304F00693
9F5FD0EFC3C50513
C5C5051300006537
04F005939E9FD0EF
A19FD0EFC0890513
494000EF27848513
0244091300842583
BDCFF0EF00090513
0009051300842583
00842703AD0FF0EF
00D7478300100513
00F706A30407E793
27848513C44FF0EF
02051E63428000EF
000065B700006437
C745859300006537
C084061306200693
975FD0EFC3C50513
C8C5051300006537
06200593969FD0EF
999FD0EFC0840513
008005133009A7F3
0181240330053573
0141248301C12083
00C1298301012903
0201011300857513
FD01011380CFC06F
000064B702912223
028124236884A783
0321202302112623
01412C2301312E23
6884849300050413
0000693702078E63
00006537000065B7
3D300693F0058593
C3C50513FA090613
000065378E1FD0EF
8D5FD0EFEB850513
FA0905133D300593
02041663905FD0EF
00040513E25FF0EF
0281240302C12083
0201290302412483
01812A0301C12983
0000806703010113
001409932B8010EF
0001262300A98433
3009397300800913
0089791300C10513
02051E632E0000EF
000065B700006A37
C245859300006537
C08A061304F00693
855FD0EFC3C50513
C5C5051300006537
04F00593849FD0EF
879FD0EFC08A0513
2F4000EF00C10513
911FF0EF0084A503
000045B70084A503
0185051300098613
1D1000EF95458593
00C105130084A703
0107E79300D74783
28C000EF00F706A3
000069B702051E63
00006537000065B7
07900693C7458593
C3C50513C0898613
00006537FD8FD0EF
FCCFD0EFC8C50513
C089851307900593
00090513FFCFD0EF
0084A783E95FB0EF
0107F79300D7C783
000064B702078E63
00006537000065B7
3F00069301858593
C3C50513FA048613
00006537F88FD0EF
F7CFD0EFEB850513
FA0485133F000593
18C010EFFACFD0EF
EA0454E340A40433
EA1FF06F00000413
00812423FF010113
FFF0079300112623
02F5126300050413
6907A503000067B7
000405135D4000EF
0081240300C12083
0000806701010113
0095051300A00413
DE9FF0EF02855533
FD9FF06F02850433
6907A503000067B7
00D5478300008067
0007986301F7F793
0015351301852503
0000051300008067
0040079300008067
00F506A300E50623
000507A300D50723
00052E2300052C23
0605202304052E23
FE01011300008067
00812C2302012303
0061202300112E23
BCDFD0EF00050413
6907A783000067B7
0687A78301C12083
0181240306F42423
0000806702010113
00812423FF010113
0005041300112623
00050663F6DFF0EF
F40FF0EF00040513
23D000EF01840513
0107E79300D44783
000067B700F406A3
028790636907A783
3005357300800513
00C1208300812403
0101011300857513
00C12083B4DFE06F
0101011300812403
0605278300008067
00812423FF010113
0005041300112623
000780E700078463
EF1FF0EF00040513
0004051302050463
00D44783EC4FF0EF
0087E79300C12083
0081240300F406A3
0000806701010113
0027F79300D44783
0004051300078663
01842783901FE0EF
01840513FC0786E3
FC1FF06F189000EF
00050E6300052503
69C7C783000067B7
40F5053300357513
0000806700A03533
0000806700100513
68878793000067B7
0087A7830147C703
0005270300E7E7B3
0005202300F71863
0000806700100513
0000806700000513
68878793000067B7
0087A7830147C703
00F5202300E7E7B3
FE01011300008067
0121282300812C23
00912A2300112E23
0005091301312623
3004347300800413
28448513000064B7
F5DFF0EF00847413
000069B702051E63
00006537000065B7
04F00693C2458593
C3C50513C0898613
00006537CD0FD0EF
CC4FD0EFC5C50513
C089851304F00593
28448513CF4FD0EF
00D94783F71FF0EF
060714630047F713
F2DFF0EF28448513
000064B702051E63
00006537000065B7
06200693C7458593
C3C50513C0848613
00006537C78FD0EF
C6CFD0EFC8C50513
C084851306200593
30042473C9CFD0EF
0181240301C12083
0101290301412483
0201011300C12983
FFB7F79300008067
0009051300F906A3
00050663D35FF0EF
910FF0EF00090513
0181240300040593
0101290301C12083
2844851300C12983
0201011301412483
FC01011384DFE06F
00068A9303512223
6886A683000066B7
02912A2302812C23
0341242303312623
0321282302112E23
0005899300050493
0441240300060A13
0000693704068E63
00006537000065B7
0509061323F00693
C3C50513F0058593
01012C2301112E23
00E1282300F12A23
00006537B90FD0EF
B84FD0EF06C50513
0509051323F00593
01C12883BB4FD0EF
0141278301812803
0401268301012703
000A061300012223
0009859300D12023
00048513000A8693
FFF00793C95FF0EF
02041A6300F40863
E11FF0EF00048513
0381240303C12083
0301290300048513
02C1298303412483
02412A8302812A03
0000806704010113
00A0061300940413
000045B702C45633
0184851395458593
4A8000EF00160613
FC010113FB9FF06F
03212823000067B7
02812C2300006937
0331262302912A23
0351222303412423
02112E2303612023
01812C2301712E23
2407849324078413
000069B724090913
00006AB700006A37
0289766300006B37
30400693094A0593
C3CA851305098613
0C4B0513A80FD0EF
30400593A78FD0EF
AA8FD0EF05098513
0004841309246463
000064B7FBCFE0EF
00006A37000069B7
FFF00B1300006AB7
00004C3700A00B93
0949859302897663
0504861332300693
A2CFD0EFC3CA0513
A24FD0EF0C4A8513
0504851332300593
07246C63A54FD0EF
03C1208303812403
0301290303412483
02812A0302C12983
02012B0302412A83
01812C0301C12B83
D51FE06F04010113
00F1222302C42783
00F1202302042783
01C4288301442783
0104270301842803
0084260300C42683
0004250300442583
00042783AFDFF0EF
030404130487AE23
02442603F0DFF06F
0004250301660863
C69FF0EF00061863
F45FF06F03040413
0376563300960613
01850513954C0593
328000EF00160613
FE010113FE1FF06F
0121282300812C23
00912A2300112E23
0005091301312623
3004347300800413
28448513000064B7
B9DFF0EF00847413
000069B702051E63
00006537000065B7
04F00693C2458593
C3C50513C0898613
00006537910FD0EF
904FD0EFC5C50513
C089851304F00593
28448513934FD0EF
00090513BB1FF0EF
000067B7A71FF0EF
032794636907A783
0181240300040593
0101290301C12083
2844851300C12983
0201011301412483
28448513D04FE06F
02051E63B41FF0EF
000065B7000064B7
C745859300006537
C084861306200693
88CFD0EFC3C50513
C8C5051300006537
06200593880FD0EF
8B0FD0EFC0848513
01C1208330042473
0141248301812403
00C1298301012903
0000806702010113
00812C23FE010113
00112E2300912A23
0005049301212823
0080041300012623
00C1051330043473
A8DFF0EF00847413
0000693702051E63
00006537000065B7
04F00693C2458593
C3C50513C0890613
00006537800FD0EF
FF5FC0EFC5C50513
C089051304F00593
00C10513824FD0EF
00C4C783AA1FF0EF
02078E630017F793
000065B700006937
1085859300006537
0E49061302900693
FB5FC0EFC3C50513
13C5051300006537
02900593FA9FC0EF
FD9FC0EF0E490513
989FF0EF00048513
68878793000067B7
069718630087A703
060794630007A783
A05FF0EF00C10513
000064B702051E63
00006537000065B7
07900693C7458593
C3C50513C0848613
00006537F51FC0EF
F45FC0EFC8C50513
C084851307900593
00040513F75FC0EF
01C12083E0CFB0EF
0141248301812403
0201011301012903
0004059300008067
B58FE0EF00C10513
000067B7FDDFF06F
000794632887A783
00000513B98FD06F
0005278300008067
0000673702050263
00E50C631F872703
0087A70300078A63
00D7073300852683
0045270300E7A423
00E7A22300F72023
0005222300052023
000067B700008067
1F478793FF010113
0007A40300812423
00F4146300112623
F89FF0EF00000413
0084278302040C63
0005546340A78533
000067B700000513
000786636987A783
0007851300A7D463
0081240300C12083
0000806701010113
FFF5451380000537
00052783FD5FF06F
02812423FD010113
01312E2302912223
0321202302112623
01512A2301412C23
0171262301612823
0005041301812423
0006049300058993
0000693702078E63
00006537000065B7
0580069317858593
C3C5051315890613
00006537DE9FC0EF
DDDFC0EFEB850513
1589051305800593
01342623E0DFC0EF
0010049300904463
3009B9F300800993
28CA051300006A37
815FF0EF0089F993
0000693702051E63
00006537000065B7
04F00693C2458593
C3C50513C0890613
00006537D89FC0EF
D7DFC0EFC5C50513
C089051304F00593
28CA0513DADFC0EF
E61FF0EF829FF0EF
000064B700950533
00A424231F44A903
00990C631F448493
00006B3700006AB7
00006C3700006BB7
0044A78302091063
00F4222300942023
0087A0230044A783
05C0006F0084A223
0207D66300892783
06100693198B0593
C3CB8513158A8613
EB8C0513D01FC0EF
06100593CF9FC0EF
D29FC0EF158A8513
0084278300892703
40F707B30AE7D863
0049278300F92423
00F4222301242023
008922230087A023
00978A630004A783
E09FF0EF00F41863
948FD0EF00000593
F34FF0EF28CA0513
0000643702051E63
00006537000065B7
06200693C7458593
C3C50513C0840613
00006537C81FC0EF
C75FC0EFC8C50513
C084051306200593
3009A9F3CA5FC0EF
0281240302C12083
0201290302412483
01812A0301C12983
01012B0301412A83
00812C0300C12B83
0000806703010113
00F4242340E787B3
EF2788E30044A783
EE5FF06F00092903
00812C23FE010113
00112E2301312623
0121282300912A23
0080041300050993
000064B730043473
0084741328C48513
02051E63E50FF0EF
000065B700006937
C245859300006537
C089061304F00693
BC5FC0EFC3C50513
C5C5051300006537
04F00593BB9FC0EF
BE9FC0EFC0890513
E64FF0EF28C48513
FEA009130009A783
0009851300078863
00000913CA5FF0EF
E14FF0EF28C48513
000064B702051E63
00006537000065B7
06200693C7458593
C3C50513C0848613
00006537B61FC0EF
B55FC0EFC8C50513
C084851306200593
30042473B85FC0EF
0181240301C12083
0141248300090513
00C1298301012903
0000806702010113
00812423FF010113
0091222300112623
0080041301212023
000064B730043473
0084741328C48513
02051E63D60FF0EF
000065B700006937
C245859300006537
C089061304F00693
AD5FC0EFC3C50513
C5C5051300006537
04F00593AC9FC0EF
AF9FC0EFC0890513
D74FF0EF28C48513
00050913C05FF0EF
D34FF0EF28C48513
000064B702051E63
00006537000065B7
06200693C7458593
C3C50513C0848613
00006537A81FC0EF
A75FC0EFC8C50513
C084851306200593
30042473AA5FC0EF
0081240300C12083
0041248300090513
0101011300012903
FE01011300008067
0121282300812C23
00112E2301412423
0131262300912A23
00058A1300050913
3004347300800413
28C48513000064B7
C74FF0EF00847413
000069B702051E63
00006537000065B7
04F00693C2458593
C3C50513C0898613
000065379E9FC0EF
9DDFC0EFC5C50513
C089851304F00593
28C48513A0DFC0EF
B19FF0EFC88FF0EF
00A7DA6300100793
000A059300A95863
E49FC0EF00090513
C34FF0EF28C48513
000064B702051E63
00006537000065B7
06200693C7458593
C3C50513C0848613
00006537981FC0EF
975FC0EFC8C50513
C084851306200593
300424739A5FC0EF
0181240301C12083
0101290301412483
00812A0300C12983
0000806702010113
02812423FD010113
0211262301412C23
0321202302912223
01512A2301312E23
0171262301612823
0191222301812423
00050A1301A12023
969FE0EF00800413
0000693730043473
0084741328C90513
02051E63B58FF0EF
000065B7000064B7
C245859300006537
C084861304F00693
8CDFC0EFC3C50513
C5C5051300006537
04F005938C1FC0EF
8F1FC0EFC0848513
28C90513000069B7
000064B7B68FF0EF
00006A372949A423
1F4A0A1328898993
00006AB726048493
00006B3700006BB7
00006CB700006C37
0009A783000A2D03
0044A5030004A683
000D0A63014D0C63
0AE7DC63008D2703
00ED242340F70733
41F7D71300D786B3
00F6B7B300A70733
00D4A02300E787B3
0009A02300F4A223
00000593985FF0EF
28C90513CC5FC0EF
02051E63AB0FF0EF
000065B7000064B7
C745859300006537
C084861306200693
FFCFC0EFC3C50513
C8C5051300006537
06200593FF0FC0EF
821FC0EFC0848513
02C1208330042473
0241248302812403
01C1298302012903
01412A8301812A03
00C12B8301012B03
00412C8300812C03
0301011300012D03
00D706B300008067
00A585B341F75593
00B6063300E6B633
000D051340E787B3
00D4A023000D2423
00F9A02300C4A223
28C9051388DFF0EF
02051663A00FF0EF
06200693C74B8593
C3CB0513C08A8613
C8CC0513F58FC0EF
06200593F50FC0EF
F80FC0EFC08A8513
00CD278330042473
00800413000D0513
30043473000780E7
0084741328C90513
02051863988FF0EF
04F00693C24C8593
C3CB0513C08A8613
00006537F08FC0EF
EFCFC0EFC5C50513
C08A851304F00593
28C90513F2CFC0EF
E6DFF06F9A8FF0EF
00912A23FE010113
00812C2300112E23
0131262301212823
3004B4F300800493
28C9051300006937
91CFF0EF0084F493
0000643702051E63
00006537000065B7
04F00693C2458593
C3C50513C0840613
00006537E90FC0EF
E84FC0EFC5C50513
C084051304F00593
28C90513EB4FC0EF
B0DFC0EF930FF0EF
26078793000067B7
0047A4030007A983
00A9B533013509B3
28C9051300850433
02051E638D8FF0EF
000065B700006937
C745859300006537
C089061306200693
E24FC0EFC3C50513
C8C5051300006537
06200593E18FC0EF
E48FC0EFC0890513
000405933004A4F3
0181240301C12083
0141248300098513
00C1298301012903
0000806702010113
2607A503000067B7
FF01011300008067
EEDFF0EF00112623
02A7B73300A00793
0101011300C12083
02A7853302B785B3
0000806700E585B3
00812C23FE010113
0000643700912A23
01212823000064B7
0141242301312623
00112E2301512223
2404849324040413
000069B700006937
00006AB700006A37
1C8985930284F663
1A89061302800693
D54FC0EFC3CA0513
D4CFC0EF0C4A8513
1A89051302800593
02946663D7CFC0EF
0181240301C12083
0101290301412483
00812A0300C12983
0000051300412A83
0000806702010113
0004051301440793
00F42C2300F42A23
01C40413BA0FB0EF
00008067F91FF06F
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
00001E1400000000
0000204000000000
0000204000000000
0000204000000000
00001D1C00000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
0000204000000000
00001C6000005F9C
00005F9C00000000
0000000000001C90
00001FB800005BFC
00005BF400000000
000061FC00002278
000055C000005F9C
0202010000000000
0404040403030303
0505050504040404
0505050505050505
0606060605050505
0606060606060606
0606060606060606
0606060606060606
0707070706060606
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0808080807070707
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0000629008080808
000062B8000062A4
000062E0000062CC
6574756D000062F4
616E796400736578
4A325B1B0063696D
4448313B35315B1B
63736544206F6D65
0A6E6F6974706972
2D2D2D2D2D2D2D2D
2D2D2D2D2D2D2D2D
6C706D69206E410A
697461746E656D65
206120666F206E6F
6E6F6974756C6F73
20656874206F7420
5020676E696E6944
68706F736F6C6968
626F72700A737265
63206128206D656C
6D2063697373616C
7268742D69746C75
636E797320646165
74617A696E6F7268
626F7270206E6F69
68540A2E296D656C
6974726170207369
6D692072616C7563
61746E656D656C70
6D6564206E6F6974
6574617274736E6F
7375206568742073
6D20666F20656761
0A656C7069746C75
6974706D65657270
20646E6120656C62
74617265706F6F63
6572687420657669
6420666F20736461
676E697265666669
7469726F69727020
0A7361202C736569
207361206C6C6577
6E61207325207325
6461657268742064
6E697065656C7320
20202020000A2E67
5652415453202020
2020202020474E49
4820202000002020
4F20474E49444C4F
204B524F4620454E
4145202000002020
205B2020474E4954
20736D2064257325
442020200000205D
4F20444550504F52
204B524F4620454E
4948542000002020
205B20474E494B4E
20736D2064257325
000000430000205D
64255B1B00000050
000000004864253B
706F736F6C696850
5B20642520726568
5D642573253A7325
4850455A00000020
2F455341425F5259
612F736F2F62696C
00632E7472657373
3A64253A73252040
747261750000000A
5F73797300000030
0000006B636F6C63
2E2E2F2E2E2F2E2E
6564756C636E692F
636F6C6E6970732F
70735F7A00682E6B
5F6B636F6C5F6E69
296C2864696C6176
4553534100000000
4146204E4F495452
205D73255B204C49
0A64253A73252040
6365520900000000
7320657669737275
0A6B636F6C6E6970
70735F7A00000000
636F6C6E755F6E69
2864696C61765F6B
746F4E090000296C
6E69707320796D20
00000A216B636F6C
425F52594850455A
686372612F455341
632F76637369722F
657268742F65726F
00000000632E6461
6F69727028282828
3D20292979746972
202626203034203D
6C64695F73695F7A
6461657268745F65
28287972746E655F
665F646165726874
7C20292929636E75
203034282828207C
203D3E202931202D
29292939322D2828
7270282820262620
2929797469726F69
322D2828203D3E20
2820262620292939
7469726F69727028
28203D3C20292979
292931202D203034
766E690900000029
6972702064696C61
252820797469726F
6F6C6C61203B2964
676E617220646577
6F74206425203A65
000000000A642520
0000238400002358
00000000000023A4
0000620400000000
0000624000006234
0000624000006240
425F52594850455A
6E72656B2F455341
6C617461662F6C65
736165720000632E
5F4B203D21206E6F
4E52454B5F525245
43494E41505F4C45
7474410900000000
7420646574706D65
65766F636572206F
61206D6F72662072
206C656E72656B20
6F632063696E6170
0A6E6F697469646E
6870657A00000000
2E312E32762D7279
35672D3337312D30
3237343531303166
202A2A2A00383034
20676E69746F6F42
4F2072796870655A
20646C6975622053
2A2A207325207325
6E69616D00000A2A
656C646900000000
4850455A00000000
2F455341425F5259
6D2F6C656E72656B
0000632E78657475
6C3E2D786574756D
6E756F635F6B636F
00005530203E2074
6574756D00000A09
72656E776F3E2D78
72656B5F203D3D20
727275632E6C656E
2E2F2E2E00746E65
72656B2F2E2E2F2E
6C636E692F6C656E
6863736B2F656475
00000000682E6465
73695F6863726121
287273695F6E695F
72656B5F00000029
727275632E6C656E
7361623E2D746E65
5F64656863732E65
212064656B636F6C
72656B5F0031203D
727275632E6C656E
7361623E2D746E65
5F64656863732E65
212064656B636F6C
656D69740030203D
30203D3E2074756F
6C6E4F0900000000
656E2D6E6F6E2079
7620657669746167
7261207365756C61
7470656363612065
000000000A2E6465
425F52594850455A
6E72656B2F455341
64656863732F6C65
657268740000632E
657361623E2D6461
5F6465646E65702E
72656B5F00006E6F
727275632E6C656E
28203D2120746E65
292A2064696F7628
695F7A2100002930
745F656C64695F73
626F5F6461657268
726874287463656A
0000000029646165
68745F73695F7A21
6174735F64616572
5F287465735F6574
632E6C656E72656B
202C746E65727275
3C3C204C55312828
0029292929342820
425F52594850455A
6E72656B2F455341
61657268742F6C65
7268540900632E64
79616D2073646165
20656220746F6E20
2064657461657263
0A73525349206E69
6572687400000000
20617461645F6461
6174735F5F203D3C
657268745F636974
5F617461645F6461
646E655F7473696C
656E750900000000
2064657463657078
646E65207473696C
6F697461636F6C20
4850455A00000A6E
2F455341425F5259
742F6C656E72656B
62615F6461657268
000000632E74726F
2D64616572687428
73752E657361623E
6F6974706F5F7265
312828202620736E
3028203C3C204C55
203D3D2029292929
7373650900005530
74206C6169746E65
6261206461657268
00000A646574726F
425F52594850455A
6E72656B2F455341
6F656D69742F6C65
00000000632E7475
6F6E645F73797321
696C5F73695F6564
6F74262864656B6E
002965646F6E3E2D
6B636974643E2D74
000030203D3E2073
425F52594850455A
6E72656B2F455341
6F706D656D2F6C65
00000000632E6C6F
5F6B5F203D3C2070
6C6F6F705F6D656D
6E655F7473696C5F
8000200000000064
000000000001C200
000061F4000014FC
02FAF080000061F4
000058A8FFFFFFF5
0000000000000000
0000000000005884
0000589C00000000
000061E400005D90
0000000000005878
0000589000000000
0000000000000000
0000624000006240
0000000000000000
0000000000000028
