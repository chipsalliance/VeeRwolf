0102829300000297
1990006F30529073
00112023FB010113
0041242300312223
0061282300512623
01C12C2300712A23
03E1202301D12E23
02A1242303F12223
02C1282302B12623
02E12C2302D12A23
0501202302F12E23
341022F305112223
300022F304512423
1F0000EF04512623
02051E6300000313
800003B7342022F3
0072F2B3FFF38393
00628A6300B00313
0000009700010513
0410006F13408093
0042829304812283
0900006F04512423
0000339700010293
0043A103B7438393
00512023FF010113
001E0E130003AE03
0003086301C3A023
03C0809300000097
342025730890006F
FFF28293800002B7
158000EF00557533
4E82829300002297
00A282B300351513
0042A3030002A503
00003317000300E7
00032383B1430313
00732023FFF38393
0002811300012283
02032E0300832383
00003297087E0863
0082A303AEC28293
0293282302832623
03332C2303232A23
0553202303432E23
0573242305632223
0593282305832623
05B32C2305A32A23
0000339702232423
0003AE0396438393
0202A30307C32623
028321030062A423
0303248302C32403
0383298303432903
04032A8303C32A03
04832B8304432B03
05032C8304C32C03
05832D8305432D03
3412907304812283
3002907304C12283
0041218300012083
00C1228300812203
0141238301012303
01C12E8301812E03
02412F8302012F03
02C1258302812503
0341268303012603
03C1278303812703
0441288304012803
3020007305010113
0000329700000073
0082A3039FC28293
0085751306C32383
00038513300522F3
0010031300008067
3442B37300A312B3
342022F300008067
0062F2B380000337
0002846300000513
0000806700150513
0200079302060063
00F04C6340C787B3
00000713FE060513
0007059300A5D533
00C5D73300008067
00F595B300C55533
FE9FF06F00B56533
0006081300058793
0005031300068893
0000273728069663
0EC5F66364470713
0CD67863000106B7
00C6B6B30FF00693
00D658B300369693
0007470301170733
0200071300D706B3
00070C6340D70733
00D556B300E797B3
00F6E5B300E61833
0108551300E51333
0108161302A5F733
0103569301065613
0107171302A5D5B3
02B607B300D766B3
00F6FE6300058713
FFF58713010686B3
00F6F6630106E863
010686B3FFE58713
02A6F7B340F686B3
0103531301031313
0107979302A6D6B3
02D605B30067E333
00B37C6300068513
FFF6851300680333
00B3746301036663
01071713FFE68513
0000059300A76733
010008B70E40006F
F3166CE301000693
F31FF06F01800693
0010069300061663
000106B702C6D833
0FF006930CD87263
008008930106F463
00D70733011856B3
0200071300074683
40D70733011686B3
410787B30A071863
0108561300100593
0108D89301081893
02C7F73301035693
0107171302C7D7B3
02F8853300D766B3
00A6FE6300078713
FFF78713010686B3
00A6F6630106E863
010686B3FFE78713
02C6F7B340A686B3
0103531301031313
0107979302C6D6B3
02D888B30067E333
01137C6300068513
FFF6851300680333
0113746301036663
01071713FFE68513
0007051300A76733
010006B700008067
F4D862E301000893
F3DFF06F01800893
00D7D5B300E81833
00D556B300E51333
00E797B301085513
00F6E8B302A5F733
0107D79301081793
02A5D5B30108D613
00C7673301071713
0005861302B786B3
0107073300D77E63
01076863FFF58613
FFE5861300D77663
40D706B301070733
0108989302A6F733
02A6D6B30108D893
02D785B301071713
00068713011767B3
010787B300B7FE63
0107E863FFF68713
FFE6871300B7F663
40B787B3010787B3
00E5E5B301061593
18D5E663EB5FF06F
04E6F46300010737
00D837330FF00813
0000283700371713
00E6D5B364480813
0005C803010585B3
00E8083302000593
02059663410585B3
EEF6ECE300100713
0015471300C53533
010005B7EEDFF06F
FCB6E0E301000713
FB9FF06F01800713
00B696B301065733
0106DE9300D766B3
03D778B30107D733
0105583300B797B3
0106979300F86333
010358130107D793
03D7573300B61633
0108E83301089893
00070E1302E78F33
00D8083301E87E63
00D86863FFF70E13
FFE70E1301E87663
41E8083300D80833
03D8583303D878B3
03078EB301089893
0107D79301031793
0008071300F8E7B3
00D787B301D7FE63
00D7E863FFF80713
FFE8071301D7F663
010E1E1300D787B3
00010EB741D787B3
FFFE881300EE6733
0107589301077333
0106561301067833
0308883303030E33
02C30333010E5693
006686B301030333
0106F46302C888B3
0106D61301D888B3
0317E663011608B3
000107B7CF179AE3
00F6F6B3FFF78793
00FE7E3301069693
01C686B300B51533
DAD57CE300000593
CC9FF06FFFF70713
0000071300000593
00002537DA5FF06F
74450513FF010113
0081242300112623
0121202300912223
00452783699000EF
0000061300100693
000005930007A783
0000041300050493
00200913000780E7
0044A783032466B3
0000059300000613
000485130047A783
000780E700140413
6D4010EF00A00513
FF010113FD9FF06F
0081242300112623
02F5046300600793
020504637B4010EF
040516637AC010EF
9FC58593000035B7
A105051300003537
2D5000EF299000EF
798010EFFFDFF06F
00003437FC051CE3
00842583C2840413
A305051300003537
00842503271000EF
FD1FF06F1B9010EF
9F858593000035B7
FB010113FB9FF06F
0491222304812423
0060079304112623
0005841300050493
000027370EA7E063
74C7071300251793
0007A78300E787B3
0000353700078067
215000EF87C50513
044427836E0010EF
00C4280301042883
0404278302F12823
0004268300442703
03C4278302F12623
0005059304842603
0384278302F12423
9005051300003537
0344278302F12223
0304278302F12023
02C4278300F12E23
0284278300F12C23
0244278300F12A23
0204278300F12823
01C4278300F12623
0184278300F12423
0144278300F12223
0084278300F12023
00040593181000EF
EA9FF0EF00048513
8A45051300003537
00003537F55FF06F
F49FF06F8C050513
0004859300003537
14D000EF8DC50513
FF010113F39FF06F
0011262300812423
3420267300050413
0016561300161613
02C7E86300500793
0026179300002737
00F707B376870713
000025370007A583
105000EF78850513
0000051300040593
000025B7EA5FF0EF
FE1FF06F78058593
00112623FF010113
00003537342025F3
0015D59300159593
0CD000EFA5850513
7A458593000025B7
E69FF0EF00400513
B3078793000037B7
00070C630007A703
0007A0230007A303
B347A503000037B7
0000806700030067
00112623FF010113
0F5000EF49D000EF
000031174F5000EF
000012B78BC10113
0051013380028293
21C0006FFD9FF0EF
01312E23FD010113
0301268300068993
0321202302812423
0006091300058413
0040061300088593
0211262302912223
00E1262300050493
0101222300F12423
00812783754010EF
00B405B3FB090593
0604A0230404AE23
02F5A823FF05F593
00C12703000027B7
8807879300412803
000017B704F5A623
0281240302C12083
0335A4239BC78793
0305AA2302E5A623
02B4A42304F5A423
0241248302012903
0301011301C12983
00C0079300008067
00C5278302F58733
00B5070300E787B3
0007A78300B75463
02E6473302000713
0027171301F67513
00F6A02300E787B3
FE01011300008067
00112E2300C10693
00C12703FBDFF0EF
00A7953300100793
01C1208300072783
00F7202300A7E7B3
0000806702010113
0085580300452783
00812423FF010113
0005041302F80833
00A4488300052503
00112623FFF00713
00E405A300912223
00C0031300000593
01F00E1301050533
0315C26302000E93
0084578300000493
00C1208306F4C463
0041248300812403
0000806701010113
00C4260302F85733
00D606B3026586B3
00C6A22300468613
00EE4E6300C6A423
0027D79300B405A3
FFC7F79300378793
FA9FF06F00158593
03D7473301F70713
0027171300A6A023
FD9FF06F00E50533
0004861300442783
02F4873300000593
0004051300042783
00E787B300148493
0047069300C42703
0087268300D7A023
0087268300D7A223
00F7242300F6A023
F51FF06FED5FF0EF
00050793FF010113
0006059300058513
0011262300068613
2FC010EF000780E7
00000513578010EF
FF01011300008067
0005041300812423
0011262304500513
0005849300912223
00048593000400E7
000400E705200513
0081240300040313
0004859300C12083
0520051300412483
0003006701010113
001787930005A783
000037B700F5A023
00030067ACC7A303
04812423FB010113
03412C2303312E23
0361282303512A23
0491222304112623
0371262305212023
0391222303812423
01B12E2303A12023
00058A9300050A13
00068B1300060993
00E0546300100413
0010079300070413
00FB146302000C13
3B9AD4B703000C13
00A00C9300100913
9FF4849300000713
00A00D1300200D93
0007146300148B93
0379D5330934F263
00190913000A8593
000A00E703050513
FFFC8C9300100713
0379F9B300100793
FCFC96E303A4D4B3
03098513000A8593
00300793000A00E7
06FB0A6341240433
0481240304C12083
0401290304412483
03812A0303C12983
03012B0303412A83
02812C0302C12B83
02012D0302412C83
0501011301C12D83
F9944CE300008067
000A8593F96DEAE3
00E12623000C0513
00190913000A00E7
F79FF06F00C12703
02000513000A8593
FFF40413000A00E7
F8DFF06FFE8048E3
04812423FB010113
0521202304912223
03412C2303312E23
0391222303512A23
01B12E2303A12023
0361282304112623
0381242303712623
0005849300050413
00068D1300060A93
FFF0091300000A13
00000C9300000993
000AC50380000DB7
04C1208304051063
0441248304812403
03C1298304012903
03412A8303812A03
02C12B8303012B03
02412C8302812C03
01C12D8302012D03
0000806705010113
02500693000C9E63
0004859336D50A63
001A8A93000400E7
06400693FA5FF06F
06A6E26310D50E63
02A6EA6303900693
0ED5746303100693
34D50A6302D00693
0CF5006303000793
02E5126302500713
0250051300048593
15C0006F000400E7
1AD50E6305800693
2EE50E6306300713
0250051300048593
00048593000400E7
FD5FF06F000AC503
16D50A6307000693
0690069302A6E063
06C006930AD50263
0680069308D50A63
FC5FF06FF6D506E3
10D5066307500693
0730071302A6EE63
000D2C03FAE518E3
000C0B93004D0B13
26051863000BC503
00F9986300300793
41790BB3418B8BB3
000B0D1327704663
078006930C80006F
07A0069312D50463
00095E63FA9FF06F
FD05091328098863
00200993F00992E3
FE0948E3EFDFF06F
02D9093300A00693
01250933FD090913
001A0A13FE1FF06F
040A1263EDDFF06F
004D0D13000D2603
0004859302065063
00C1202302D00513
00012603000400E7
40C00633FFF90913
0009869300090713
0004051300048593
03C0006FCA1FF0EF
FAEA0EE300100713
FF87F713007D0793
0047268300072603
01B6073300870D13
00D7073300C73733
00048593FA0700E3
C01FF0EF00040513
E59FF06F00000C93
000D2603000A1863
F9DFF06F004D0D13
FEEA08E300100713
FF87F713007D0793
0007260300870D13
FC0710E300472703
FFF7C793800007B7
FB1FF06FF6C7F8E3
0300051300048593
00048593000400E7
000400E707800513
0010099300800913
0B46C26300100693
00012423000D2783
00F12223004D0D13
00000B9301000C13
0100089300012023
0081258300412503
002B1613FFF88B13
9CCFF0EF01112623
0805186300F57513
0300069300012783
00C1288300079863
08F8966300100793
0185151300A68533
4185551300048593
001B8B93000400E7
00300693040B1863
D6D998E300000C93
41770BB300191713
00048593F17054E3
000400E702000513
FEDFF06FFFFB8B93
FF87F693007D0793
00868D130006A783
0046A78300F12223
F55FF06F00F12423
000B089301912023
00900793F59FF06F
F8A7E2E305700693
F7DFF06F03000693
00F12623FFFC0793
0010079301894C63
0004859300F99C63
000400E703000513
FC1FF06F00C12C03
FEF99AE300200793
0200051300048593
00048593FE5FF06F
000400E7001B8B93
00048593D81FF06F
000400E702000513
D85FF06FFFFB8B93
00048593000D2503
000400E7004D0B13
00000A13D75FF06F
00000993FFF00913
C89FF06F00100C93
C81FF06F00300993
C79FF06F00100993
00050613FE010113
0005869300001537
00C10593C5050513
0001262300112E23
01C12083BA1FF0EF
0000806702010113
02B12223FC010113
00112E2302410593
02D1262302C12423
02F12A2302E12823
03112E2303012C23
FA5FF0EF00B12623
0401011301C12083
0000806700008067
3007A7F300800793
0000806710500073
00A7953300100793
0000806730452573
00A7953300100793
0000806730453573
3007B7F300800793
3440507330405073
FF01011300008067
0011262300700513
800016B7FD1FF0EF
0003D7370186A783
00E787B309070713
00F6AC2300700513
00C12083FA1FF0EF
0101011300100513
FF01011314C0106F
0011262300700513
800016B7F91FF0EF
0003D7370186A783
00E787B309070713
00F6AC2300700513
00C12083F61FF0EF
0101011300000513
0000806700008067
0000806700000513
0005C70300054783
0007966300E79463
0000806740E78533
0015859300150513
0FF5F693FE1FF06F
0037F71300050793
0FF5F59304071863
00B765B300859713
00B765B301059713
0007871300C78333
40E308B300300813
0026571303186E63
00B787B300271593
02B70733FFC00593
00E7873300C70733
0000806702E79463
00178793FE060EE3
FFF60613FED78FA3
00470713F9DFF06F
FB9FF06FFEB72E23
FED78FA300178793
00852703FD1FF06F
00B7E5B30026F793
04059A6300072503
00C7963300100793
FEA0051300452783
0407806300F677B3
FDD00513F7E6F793
0806F51302079A63
00050A6300472783
00C7222300F66633
0000806700000513
00F67633FFF64613
0000806700C72223
00008067FDD00513
0007A50300852783
000528830047A783
0205906300452803
00C7173300100713
FEA0051300E87833
0006846302080C63
0080071300080693
0008A60330073773
00F647B300877713
0107F7B300D7C7B3
00F8A02300C7C7B3
0000051330072773
0085250300008067
0045250300052703
0007A78300072783
0047250300A7C7B3
0205986300A7F7B3
0017F79300C7D7B3
0010079300F6A023
0047260300C797B3
0007946300C7F7B3
00058513FEA00593
00F6A02300008067
FF1FF06F00000593
0085278300052703
00E7A02300872703
A8C78793000037B7
0000051300F52223
0025171300008067
00150513000037B7
00251513AA878793
00E78733FF010113
0081242300A787B3
0007240300912223
001126230007A483
00C1208300946C63
0041248300812403
0000806701010113
0004051300042783
000780E70047A783
0004222300050463
FCDFF06F00C40413
000037B7FF010113
000034B700912223
0011262300812423
01212023AE878413
B0C48493AE878793
0005091300941C63
0294146300078413
0440006F00000413
0007086300442703
0007270300042703
00C4041302A70863
00442783FD1FF06F
00C4041300079663
00042783FCDFF06F
0007A58300090513
FE0514E3D21FF0EF
00C1208300040513
0041248300812403
0101011300012903
0000353700008067
B2050613000037B7
40C78633C5478793
B205051300000593
FF010113D05FF06F
0011262300200513
00300513ECDFF0EF
201000EFEC5FF0EF
000037B7874FF0EF
00C7C703BB878793
00E78623FFE77713
0101011300C12083
F601011300008067
000047B708812C23
0931262300003437
C2840993A6078793
0101079300F9A223
0000059307000613
08112E2300078513
0921282308912A23
00100713C85FF0EF
0000051300A9A423
E49FF0EF00E10EA3
E41FF0EF00100513
00F11E2310100793
000037B7638000EF
00003937ABC78793
000016B700F12223
000035B700100793
00F12023BB890493
0000079300000713
0000081300000893
4000061365468693
BB890513C6058593
079000EF0299A023
C284041300D4C783
00E486A3FFB7F713
00079A6301B7F793
000796630184A783
2DC000EFBB890513
AC478793000037B7
0000353700F12223
000026B700100793
B4850493000035B7
00F0089300F12023
0000079300000813
5546869300000713
0605859320000613
009000EFB4850513
0094262300D4C783
FFB7F79300800513
000037B700F486A3
00F42C23C4078793
3005357300F42E23
A45FE0EF00857513
0005278300452703
00E7A22300F72023
0005222300052023
00D5478300008067
0007986301F7F793
0015351301852503
0000051300008067
FF01011300008067
AFDFF0EF00112623
B3C7A783000037B7
0000373700C12083
C2A72C2300A78533
0007851300000593
3810006F01010113
00812423FF010113
0080041300112623
000037B730043473
00950513C207AC23
02F5453300A00793
00847413000037B7
000037B7B2A7AE23
F91FF0EFB2B7AC23
00C1208330042473
0101011300812403
FF01011300008067
0091222300812423
0005049300112623
3004347300800413
00D4C783F21FF0EF
FFD7F79300847413
3004247300F486A3
0081240300C12083
004124830004A423
0000806701010113
C287A783000037B7
0005851300079663
0085F593921FE06F
000080673005A5F3
C287270300003737
905FE06F00071463
3007A7F300857793
0080051300008067
0085751330053573
00800793FD9FF06F
000037373007B7F3
00F6C703C3072683
00E687A3FFF70713
3007A7F30087F793
0005278300008067
0000079300F51463
0000806700078513
00812C23FE010113
00912A2300003437
C284051300050493
00112E2302450513
C2840413FCDFF0EF
00C4250300051463
02049A6300842783
01F7771300D7C703
00E7D68302071463
00D77E6307F00713
01C1208302F42023
0141248301812403
0000806702010113
00A1262300F50863
00C12503E35FF0EF
FD9FF06F02A42023
00812423FF010113
0080041300112623
000037B730043473
00100513C307A703
00F7478300847413
00F707A300178793
30042473F51FF0EF
00C1208300812403
EF1FF06F01010113
00812423FF010113
0080041300112623
0000373730043473
0247A783C2870793
C4C68693000036B7
C287071300847413
04078E6306D78063
00E5060302872583
0506506300E78803
00F520230047A703
00A7202300E52223
00D5478300A7A223
00F506A30407E793
ECDFF0EF00000513
00C1208330042473
0101011300812403
00B7866300008067
FA079AE30007A783
00D5202302872783
0287278300F52223
02A7242300A7A023
FF052783FB5FF06F
00812423FF010113
0011262301212023
0005041300912223
02078663FE850913
3004B4F300800493
CC5FF0EF00090513
0084F493FF544783
FEF40AA3FFD7F793
FE0428233004A4F3
00090513FF544783
FEF40AA3FEB7F793
02050063CB5FF0EF
00C1208300812403
0009051300412483
0101011300012903
00C12083ED9FF06F
0041248300812403
0101011300012903
FF01011300008067
0091222300812423
0005041300112623
3004B4F300800493
00003737C41FF0EF
0247A783C2870793
C4C68693000036B7
C28707130084F493
0607846306D78663
00E4060302872583
04A6566300E78503
00F420230047A683
0086A02300D42223
00D447830087A223
0407E79300872503
00F406A340850533
D75FF0EF00153513
00C120833004A4F3
0041248300812403
0000806701010113
0007A78300B78663
02872783FA0794E3
00F4222300D42023
0087A02302872783
FA9FF06F02872423
B3C7A783000037B7
000037B706078663
0087A703C2878793
00E7560307F00693
000036B704C6EA63
B386A68300E70603
000036B704D64263
02D70C63AE46A683
0206986301872683
02D540630107A683
00070513FF010113
EE1FF0EF00112623
0101011300C12083
40A686B3B6DFF06F
0000806700D7A823
00812423FF010113
0011262300912223
0080041300050493
00D5478330043473
0407F79300847413
AF5FF0EF00078A63
FBF7F79300D4C783
000037B700F486A3
40950533C307A503
C6DFF0EF00153513
00C1208330042473
0041248300812403
0000806701010113
C2878793000037B7
02E7A22302478713
0000059302E7A423
B0DFF06F00000513
00812423FF010113
C284079300003437
000037B70087A703
00112623AE47A783
06F7026300912223
00800493C2840413
008425033004B4F3
A5DFF0EF0084F493
000036B702442783
00842703C4C68693
0607806306D78263
00E7058302842603
04A5D26300E78503
00F720230047A683
00E6A02300D72223
0010051300E7A223
3004A4F3BB1FF0EF
3005357300800513
00C1208300812403
0085751300412483
C34FE06F01010113
0007A78300F60663
02842783FA0798E3
00F7222300D72023
00E7A02302842783
FB1FF06F02E42423
02112623FD010113
0291222302812423
01312E2303212023
00A1262302051663
00C12503F11FF0EF
0281240302C12083
0201290302412483
0301011301C12983
0095041300008067
02A4443300A00513
008009936D8000EF
00A404B300140413
000039373009B9F3
00892503C2890913
00892503E39FF0EF
00040613000025B7
01850513AF458593
008927033D8000EF
00D747830089F513
00F706A30107E793
684000EFB68FE0EF
0000051340A484B3
3E800513F6905CE3
0640061302A495B3
02A4853300000693
F5DFF06FBC8FE0EF
C307A503000037B7
00D5478300008067
0007986301F7F793
0015351301852503
0000051300008067
000037B700008067
00A03533C287A503
000037B700008067
00C7C503C307A783
0000806700157513
00812423FF010113
0091222300112623
3004347300800413
0084741300D54783
00071E630047F713
00C1208330042473
0041248300812403
0000806701010113
00F506A3FFB7F793
F71FF0EF00050493
0004851300050663
00040593AB1FF0EF
00C1208300812403
0000353700412483
01010113C5450513
FE010113941FF06F
00812C2302012303
0061202300112E23
9EDFE0EF00050413
C307A783000037B7
0687A78301C12083
0181240306F42423
0000806702010113
FF01011306052783
0011262300812423
0007846300050413
00040513000780E7
02050463EE5FF0EF
CA5FF0EF00040513
00C1208300D44783
00F406A30087E793
0101011300812403
00D4478300008067
000786630027F793
859FF0EF00040513
FC0786E301842783
2FC000EF01840513
FD010113FC1FF06F
03212023000037B7
0281242300003937
0211262302912223
01412C2301312E23
B0C78493B0C78413
03246E63B0C90913
8A1FF0EF00048413
00A00993FFF00493
0724646300002A37
02C1208302812403
0201290302412483
01812A0301C12983
92DFF06F03010113
00F1222302C42783
00F1202302042783
01C4288301442783
0104270301842803
0084260300C42683
0004250300442583
00042783EB5FF0EF
030404130487AE23
02442603F85FF06F
0004250300960863
E15FF0EF00061863
F81FF06F03040413
0336463300960613
01850513AF4A0593
134000EF00160613
00D50623FE1FF06F
00B5072300C506A3
00052C23000507A3
0000806700052E23
02112623FD010113
3005B5F300800593
00B126230085F593
00C12583E71FF0EF
F64FF0EF01C10513
0301011302C12083
000037B700008067
00079463B407A783
00000513978FF06F
0005278300008067
0000373702050263
00E50C63AD472703
0087A70300078A63
00D7073300852683
0045270300E7A423
00E7A22300F72023
0005222300052023
000037B700008067
FF010113B447C783
0081242300112623
FFF0051300912223
8000053700079663
000037B7FFF54513
0007A403AD078793
0204026302F40463
F69FF0EF00842483
0000051340A484B3
008424030004C863
40A40533F55FF0EF
C387A783000037B7
00A7D46300078663
00C1208300078513
0041248300812403
0000806701010113
00812C23FE010113
00112E2300912A23
00C1262300050413
0080049300B52623
F01FF0EF3004B4F3
0084F49300C12603
0010061300C04463
AD07A703000037B7
00C4242300A60633
00F70663AD078793
020710630047A583
00F420230047A703
0047A70300E42223
0087A22300872023
0087260302C0006F
04C6D86300842683
00D7242340D606B3
00E4202300472683
0086A02300D42223
0007A70300872223
00E4186300F70A63
00000593ED5FF0EF
3004A4F3FF5FE0EF
0181240301C12083
0201011301412483
40C686B300008067
F8B702E300D42423
F79FF06F00072703
00812423FF010113
0080041300112623
0005278330043473
0207806300847413
00000513E3DFF0EF
00C1208330042473
0101011300812403
FEA0051300008067
FF010113FE9FF06F
0081242300112623
3007B47300800793
00847793E45FF0EF
00C120833007A7F3
0101011300812403
FE01011300008067
00912A2300812C23
0005049300112E23
0080041300B12623
E09FF0EF30043473
00C1258300847413
0010079300A4DA63
0004851300A7D663
30042473F15FE0EF
0181240301C12083
0201011301412483
FE01011300008067
00912A2300812C23
0121282300112E23
0141242301312623
0005049301512223
FFCFF0EF00800413
000039B730043473
0000393700003A37
00847413B499A023
AD0A0A13B4098993
00800A93B2090913
0009A783000A2483
0049250300092683
00048A6301448C63
06E7D0630084A703
00E4A42340F70733
41F7D71300D786B3
00F6B7B300A70733
00D9202300E787B3
0009A02300F92223
00000593D35FF0EF
30042473E55FE0EF
0181240301C12083
0101290301412483
00812A0300C12983
0201011300412A83
00D706B300008067
00A585B341F75593
00B6063300E6B633
0004A42340E787B3
00D9202300048513
00F9A02300C92223
30042473C95FF0EF
0004851300C4A783
300AB473000780E7
F3DFF06F00847413
B207A503000037B7
FF01011300008067
0011262300812423
300437F300800413
00A04463E3DFF0EF
0010059300100513
CE5FE0EFE5DFF0EF
FF010113FE5FF06F
0091222300812423
000034B700003437
B0C4041300112623
00946E63B0C48493
0081240300C12083
0000051300412483
0000806701010113
0004051301440793
00F42C2300F42A23
01C40413D08FE0EF
00008067FCDFF06F
0000093800000000
0000093800000000
0000093800000000
0000093800000000
0000093800000000
0000093800000000
0000093800000000
000012A400000000
0000150800002744
00002A8000002AD8
00000000000012E4
00002584000027A0
0202010000000000
0404040403030303
0505050504040404
0505050505050505
0606060605050505
0606060606060606
0606060606060606
0606060606060606
0707070706060606
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0707070707070707
0808080807070707
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
0808080808080808
3044454C08080808
0000081000000000
000008C8000008C8
0000081000000804
000008BC000008B0
00002814000027F4
0000284400002830
0000286800002850
006E776F6E6B6E75
6F69747065637845
206573756163206E
0A29642528207325
DEADBAAD00000000
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
DEADBAADDEADBAAD
74736E49DEADBAAD
206E6F6974637572
2073736572646461
6E67696C6173696D
74736E4900006465
206E6F6974637572
6620737365636341
00000000746C7561
206C6167656C6C49
7463757274736E69
61657242006E6F69
0000746E696F706B
6464612064616F4C
73696D2073736572
0064656E67696C61
6363612064616F4C
6C75616620737365
2A2A2A2A00000074
206C656E72654B20
697461636F6C6C41
756C696146206E6F
2A2A2A2A20216572
2A2A2A2A0000000A
6C656E72654B202A
2A202153504F4F20
0000000A2A2A2A2A
654B202A2A2A2A2A
6E6150206C656E72
2A2A2A2A20216369
2A2A2A2A00000A2A
6E776F6E6B6E5520
45206C6174614620
21642520726F7272
00000A2A2A2A2A20
20746E6572727543
4920646165726874
460A7025203D2044
20676E69746C7561
7463757274736E69
72646461206E6F69
7830203D20737365
3A617220200A7825
6720207825783020
2078257830203A70
257830203A707420
30203A3074202078
317420200A782578
202078257830203A
78257830203A3274
7830203A33742020
203A347420207825
7420200A78257830
2078257830203A35
257830203A367420
30203A3061202078
3A31612020782578
20200A7825783020
78257830203A3261
7830203A33612020
203A346120207825
3561202078257830
200A78257830203A
257830203A366120
30203A3761202078
000000000A782578
6573736500525349
6874206C6169746E
0000000064616572
6166206C61746146
25206E6920746C75
6E6E697053202173
000A2E2E2E676E69
6166206C61746146
74206E6920746C75
7025206461657268
6974726F62412021
000000000A2E676E
73756F6972757053
75727265746E6920
6365746564207470
5152492021646574
0000000A6425203A
636F6C635F737973
000013DC0000006B
000014AC00001448
0000000000000000
0000000000000000
00002B0000002AE8
00002B0C00002B0C
6E69616D00002B0C
656C646900000000
00000BFCFFFFFF00
00002AD000002AD0
0000000180001010
00002B48FFFFFFF5
0000000000002638
0000262000000000
00002B2800000000
000000000000262C
00002B0C00000000
0000000000002B0C
0000000F00000000
