08000E1380002537
01B00E9301C50623
00300E1301D50023
08700E1301C50623
0005022301C50423
0005828306000593
0015859301C000EF
FE029AE300058283
800015B70000006F
01450F8300958593
FE0F8CE3020FFF93
0000806700550023
7375462B52656556
636F7220436F5365
00000000000A736B
