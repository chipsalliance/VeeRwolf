0105051380001537
0055002300100337
000073B30012C293
FE731EE300138393
00000000FEDFF06F
